
module conv_16_4_16_1 ( clk, reset, s_data_in_x, s_valid_x, s_ready_x, 
        m_data_out_y, m_valid_y, m_ready_y );
  input [15:0] s_data_in_x;
  output [15:0] m_data_out_y;
  input clk, reset, s_valid_x, m_ready_y;
  output s_ready_x, m_valid_y;
  wire   w_conv_done, e_acc, c_acc, \mx/N29 , \mx/N28 , \mx/N26 , \mx/N25 ,
         \mx/N24 , \mx/N21 , \mx/N19 , \mx/N18 , \mx/N17 , \mx/N16 , \mx/N15 ,
         \mx/N14 , \mx/mem[15][15] , \mx/mem[15][14] , \mx/mem[15][13] ,
         \mx/mem[15][12] , \mx/mem[15][11] , \mx/mem[15][10] , \mx/mem[15][9] ,
         \mx/mem[15][8] , \mx/mem[15][7] , \mx/mem[15][6] , \mx/mem[15][5] ,
         \mx/mem[15][4] , \mx/mem[15][3] , \mx/mem[15][2] , \mx/mem[15][1] ,
         \mx/mem[15][0] , \mx/mem[14][15] , \mx/mem[14][14] , \mx/mem[14][13] ,
         \mx/mem[14][12] , \mx/mem[14][11] , \mx/mem[14][10] , \mx/mem[14][9] ,
         \mx/mem[14][8] , \mx/mem[14][7] , \mx/mem[14][6] , \mx/mem[14][5] ,
         \mx/mem[14][4] , \mx/mem[14][3] , \mx/mem[14][2] , \mx/mem[14][1] ,
         \mx/mem[14][0] , \mx/mem[13][15] , \mx/mem[13][14] , \mx/mem[13][13] ,
         \mx/mem[13][12] , \mx/mem[13][11] , \mx/mem[13][10] , \mx/mem[13][9] ,
         \mx/mem[13][8] , \mx/mem[13][7] , \mx/mem[13][6] , \mx/mem[13][5] ,
         \mx/mem[13][4] , \mx/mem[13][3] , \mx/mem[13][2] , \mx/mem[13][1] ,
         \mx/mem[13][0] , \mx/mem[12][15] , \mx/mem[12][14] , \mx/mem[12][13] ,
         \mx/mem[12][12] , \mx/mem[12][11] , \mx/mem[12][10] , \mx/mem[12][9] ,
         \mx/mem[12][8] , \mx/mem[12][7] , \mx/mem[12][6] , \mx/mem[12][5] ,
         \mx/mem[12][4] , \mx/mem[12][3] , \mx/mem[12][2] , \mx/mem[12][1] ,
         \mx/mem[12][0] , \mx/mem[11][15] , \mx/mem[11][14] , \mx/mem[11][13] ,
         \mx/mem[11][12] , \mx/mem[11][11] , \mx/mem[11][10] , \mx/mem[11][9] ,
         \mx/mem[11][8] , \mx/mem[11][7] , \mx/mem[11][6] , \mx/mem[11][5] ,
         \mx/mem[11][4] , \mx/mem[11][3] , \mx/mem[11][2] , \mx/mem[11][1] ,
         \mx/mem[11][0] , \mx/mem[10][15] , \mx/mem[10][14] , \mx/mem[10][13] ,
         \mx/mem[10][12] , \mx/mem[10][11] , \mx/mem[10][10] , \mx/mem[10][9] ,
         \mx/mem[10][8] , \mx/mem[10][7] , \mx/mem[10][6] , \mx/mem[10][5] ,
         \mx/mem[10][4] , \mx/mem[10][3] , \mx/mem[10][2] , \mx/mem[10][1] ,
         \mx/mem[10][0] , \mx/mem[9][15] , \mx/mem[9][14] , \mx/mem[9][13] ,
         \mx/mem[9][12] , \mx/mem[9][11] , \mx/mem[9][10] , \mx/mem[9][9] ,
         \mx/mem[9][8] , \mx/mem[9][7] , \mx/mem[9][6] , \mx/mem[9][5] ,
         \mx/mem[9][4] , \mx/mem[9][3] , \mx/mem[9][2] , \mx/mem[9][1] ,
         \mx/mem[9][0] , \mx/mem[8][15] , \mx/mem[8][14] , \mx/mem[8][13] ,
         \mx/mem[8][12] , \mx/mem[8][11] , \mx/mem[8][10] , \mx/mem[8][9] ,
         \mx/mem[8][8] , \mx/mem[8][7] , \mx/mem[8][6] , \mx/mem[8][5] ,
         \mx/mem[8][4] , \mx/mem[8][3] , \mx/mem[8][2] , \mx/mem[8][1] ,
         \mx/mem[8][0] , \mx/mem[7][15] , \mx/mem[7][14] , \mx/mem[7][13] ,
         \mx/mem[7][12] , \mx/mem[7][11] , \mx/mem[7][10] , \mx/mem[7][9] ,
         \mx/mem[7][8] , \mx/mem[7][7] , \mx/mem[7][6] , \mx/mem[7][5] ,
         \mx/mem[7][4] , \mx/mem[7][3] , \mx/mem[7][2] , \mx/mem[7][1] ,
         \mx/mem[7][0] , \mx/mem[6][15] , \mx/mem[6][14] , \mx/mem[6][13] ,
         \mx/mem[6][12] , \mx/mem[6][11] , \mx/mem[6][10] , \mx/mem[6][9] ,
         \mx/mem[6][8] , \mx/mem[6][7] , \mx/mem[6][6] , \mx/mem[6][5] ,
         \mx/mem[6][4] , \mx/mem[6][3] , \mx/mem[6][2] , \mx/mem[6][1] ,
         \mx/mem[6][0] , \mx/mem[5][15] , \mx/mem[5][14] , \mx/mem[5][13] ,
         \mx/mem[5][12] , \mx/mem[5][11] , \mx/mem[5][10] , \mx/mem[5][9] ,
         \mx/mem[5][8] , \mx/mem[5][7] , \mx/mem[5][6] , \mx/mem[5][5] ,
         \mx/mem[5][4] , \mx/mem[5][3] , \mx/mem[5][2] , \mx/mem[5][1] ,
         \mx/mem[5][0] , \mx/mem[4][15] , \mx/mem[4][14] , \mx/mem[4][13] ,
         \mx/mem[4][12] , \mx/mem[4][11] , \mx/mem[4][10] , \mx/mem[4][9] ,
         \mx/mem[4][8] , \mx/mem[4][7] , \mx/mem[4][6] , \mx/mem[4][5] ,
         \mx/mem[4][4] , \mx/mem[4][3] , \mx/mem[4][2] , \mx/mem[4][1] ,
         \mx/mem[4][0] , \mx/mem[3][15] , \mx/mem[3][14] , \mx/mem[3][13] ,
         \mx/mem[3][12] , \mx/mem[3][11] , \mx/mem[3][10] , \mx/mem[3][9] ,
         \mx/mem[3][8] , \mx/mem[3][7] , \mx/mem[3][6] , \mx/mem[3][5] ,
         \mx/mem[3][4] , \mx/mem[3][3] , \mx/mem[3][2] , \mx/mem[3][1] ,
         \mx/mem[3][0] , \mx/mem[2][15] , \mx/mem[2][14] , \mx/mem[2][13] ,
         \mx/mem[2][12] , \mx/mem[2][11] , \mx/mem[2][10] , \mx/mem[2][9] ,
         \mx/mem[2][8] , \mx/mem[2][7] , \mx/mem[2][6] , \mx/mem[2][5] ,
         \mx/mem[2][4] , \mx/mem[2][3] , \mx/mem[2][2] , \mx/mem[2][1] ,
         \mx/mem[2][0] , \mx/mem[1][15] , \mx/mem[1][14] , \mx/mem[1][13] ,
         \mx/mem[1][12] , \mx/mem[1][11] , \mx/mem[1][10] , \mx/mem[1][9] ,
         \mx/mem[1][8] , \mx/mem[1][7] , \mx/mem[1][6] , \mx/mem[1][5] ,
         \mx/mem[1][4] , \mx/mem[1][3] , \mx/mem[1][2] , \mx/mem[1][1] ,
         \mx/mem[1][0] , \mx/mem[0][15] , \mx/mem[0][14] , \mx/mem[0][13] ,
         \mx/mem[0][12] , \mx/mem[0][11] , \mx/mem[0][10] , \mx/mem[0][9] ,
         \mx/mem[0][8] , \mx/mem[0][7] , \mx/mem[0][6] , \mx/mem[0][5] ,
         \mx/mem[0][4] , \mx/mem[0][3] , \mx/mem[0][2] , \mx/mem[0][1] ,
         \mx/mem[0][0] , \mf/N17 , \mf/N15 , \mf/N14 , \mf/N13 , \mf/N12 ,
         \cx/overflow , \cc/N56 , \cc/hold_state , \cc/en_val_y , \conv/N146 ,
         \conv/N145 , \conv/N144 , \conv/N143 , \conv/N142 , \conv/N141 ,
         \conv/N140 , \conv/N139 , \conv/N138 , \conv/N137 , \conv/N136 ,
         \conv/N135 , \conv/N134 , \conv/N133 , \conv/N132 , \conv/N125 ,
         \conv/N124 , \conv/N123 , \conv/N122 , \conv/N121 , \conv/N120 ,
         \conv/N119 , \conv/N118 , \conv/N117 , \conv/N116 , \conv/N115 ,
         \conv/N114 , \conv/N113 , \conv/N112 , \conv/N111 , \conv/N110 , n654,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n923, n924, n925, n926, n927, n928, n929, \DP_OP_65J1_123_5677/n1047 ,
         \DP_OP_65J1_123_5677/n1044 , n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378;
  wire   [3:0] w_write_addr_x;
  wire   [3:0] w_read_addr_x;
  wire   [1:0] w_read_addr_f;
  wire   [15:0] w_to_multx;
  wire   [15:0] w_to_multf;
  wire   [3:0] \cc/number_x ;
  wire   [15:0] \conv/prev_output ;
  assign m_data_out_y[15] = 1'b0;

  DFF_X1 \mx/data_out_reg[4]  ( .D(\mx/N25 ), .CK(clk), .Q(w_to_multx[4]) );
  DFF_X1 \mx/data_out_reg[8]  ( .D(\mx/N21 ), .CK(clk), .Q(w_to_multx[8]), 
        .QN(n1021) );
  DFF_X1 \mx/data_out_reg[10]  ( .D(\mx/N19 ), .CK(clk), .Q(w_to_multx[10]), 
        .QN(n1022) );
  DFF_X1 \mx/data_out_reg[12]  ( .D(\mx/N17 ), .CK(clk), .Q(w_to_multx[12]), 
        .QN(n995) );
  DFF_X1 \mx/data_out_reg[14]  ( .D(\mx/N15 ), .CK(clk), .Q(w_to_multx[14]), 
        .QN(n992) );
  DFF_X1 \mx/data_out_reg[15]  ( .D(\mx/N14 ), .CK(clk), .Q(w_to_multx[15]), 
        .QN(n1013) );
  DFF_X1 \mf/z_reg[5]  ( .D(\mf/N15 ), .CK(clk), .Q(w_to_multf[5]), .QN(n946)
         );
  DFF_X1 \cc/m_addr_read_f_reg[0]  ( .D(n920), .CK(clk), .Q(w_read_addr_f[0])
         );
  DFF_X1 \cc/en_val_y_reg  ( .D(n929), .CK(clk), .Q(\cc/en_val_y ) );
  DFF_X1 \cc/en_acc_reg  ( .D(\cc/N56 ), .CK(clk), .Q(e_acc) );
  DFF_X1 \cc/conv_done_reg  ( .D(n926), .CK(clk), .Q(w_conv_done) );
  DFF_X1 \cc/number_x_reg[2]  ( .D(n916), .CK(clk), .Q(\cc/number_x [2]) );
  DFF_X1 \cc/m_addr_read_x_reg[3]  ( .D(n911), .CK(clk), .Q(w_read_addr_x[3])
         );
  DFF_X1 \conv/prev_output_reg[11]  ( .D(\conv/N121 ), .CK(clk), .QN(n2100) );
  DFF_X1 \cc/hold_state_reg  ( .D(n654), .CK(clk), .Q(\cc/hold_state ) );
  DFF_X1 \mx/data_out_reg[1]  ( .D(\mx/N28 ), .CK(clk), .Q(
        \DP_OP_65J1_123_5677/n1047 ), .QN(n1039) );
  DFF_X1 \mx/data_out_reg[5]  ( .D(\mx/N24 ), .CK(clk), .Q(w_to_multx[5]), 
        .QN(n1018) );
  DFF_X1 \conv/m_data_out_y_reg[9]  ( .D(\conv/N141 ), .CK(clk), .Q(
        m_data_out_y[9]) );
  DFF_X1 \mx/data_out_reg[9]  ( .D(n1038), .CK(clk), .Q(n2104), .QN(
        w_to_multx[9]) );
  DFF_X1 \mx/data_out_reg[7]  ( .D(n1037), .CK(clk), .Q(n2378), .QN(
        \DP_OP_65J1_123_5677/n1044 ) );
  DFF_X1 \mf/z_reg[15]  ( .D(\mf/N17 ), .CK(clk), .Q(w_to_multf[7]), .QN(
        w_to_multf[15]) );
  DFF_X1 \mx/data_out_reg[6]  ( .D(n1036), .CK(clk), .Q(n2106), .QN(
        w_to_multx[6]) );
  DFF_X1 \conv/m_data_out_y_reg[7]  ( .D(\conv/N139 ), .CK(clk), .Q(
        m_data_out_y[7]) );
  DFF_X1 \conv/m_data_out_y_reg[13]  ( .D(\conv/N145 ), .CK(clk), .Q(
        m_data_out_y[13]) );
  DFF_X1 \cc/clr_acc_reg  ( .D(n928), .CK(clk), .Q(c_acc), .QN(n2111) );
  DFF_X1 \cc/m_valid_y_reg  ( .D(n927), .CK(clk), .Q(m_valid_y), .QN(n2114) );
  DFF_X1 \cx/m_addr_x_reg[0]  ( .D(n923), .CK(clk), .Q(w_write_addr_x[0]), 
        .QN(n2108) );
  DFF_X1 \cc/number_x_reg[0]  ( .D(n918), .CK(clk), .Q(\cc/number_x [0]), .QN(
        n2115) );
  DFF_X1 \cx/overflow_reg  ( .D(n924), .CK(clk), .Q(\cx/overflow ), .QN(n2110)
         );
  DFF_X1 \cc/number_x_reg[1]  ( .D(n917), .CK(clk), .Q(\cc/number_x [1]), .QN(
        n2118) );
  DFF_X1 \cc/m_addr_read_f_reg[1]  ( .D(n919), .CK(clk), .Q(w_read_addr_f[1]), 
        .QN(n2117) );
  DFF_X1 \cx/m_addr_x_reg[1]  ( .D(n2121), .CK(clk), .Q(n2107), .QN(
        w_write_addr_x[1]) );
  DFF_X1 \cx/m_addr_x_reg[2]  ( .D(n921), .CK(clk), .Q(w_write_addr_x[2]), 
        .QN(n2112) );
  DFF_X1 \cc/number_x_reg[3]  ( .D(n915), .CK(clk), .Q(\cc/number_x [3]), .QN(
        n2120) );
  DFF_X1 \cx/m_addr_x_reg[3]  ( .D(n925), .CK(clk), .Q(w_write_addr_x[3]), 
        .QN(n2109) );
  DFF_X1 \cc/m_addr_read_x_reg[0]  ( .D(n914), .CK(clk), .Q(w_read_addr_x[0]), 
        .QN(n2113) );
  DFF_X1 \cc/m_addr_read_x_reg[1]  ( .D(n913), .CK(clk), .Q(w_read_addr_x[1]), 
        .QN(n2116) );
  DFF_X1 \cc/m_addr_read_x_reg[2]  ( .D(n912), .CK(clk), .Q(w_read_addr_x[2]), 
        .QN(n2119) );
  DFF_X1 \mx/mem_reg[6][15]  ( .D(n2233), .CK(clk), .QN(\mx/mem[6][15] ) );
  DFF_X1 \mx/mem_reg[6][14]  ( .D(n2232), .CK(clk), .QN(\mx/mem[6][14] ) );
  DFF_X1 \mx/mem_reg[6][13]  ( .D(n2231), .CK(clk), .QN(\mx/mem[6][13] ) );
  DFF_X1 \mx/mem_reg[6][12]  ( .D(n2230), .CK(clk), .QN(\mx/mem[6][12] ) );
  DFF_X1 \mx/mem_reg[6][11]  ( .D(n2229), .CK(clk), .QN(\mx/mem[6][11] ) );
  DFF_X1 \mx/mem_reg[6][10]  ( .D(n2228), .CK(clk), .QN(\mx/mem[6][10] ) );
  DFF_X1 \mx/mem_reg[6][9]  ( .D(n2227), .CK(clk), .QN(\mx/mem[6][9] ) );
  DFF_X1 \mx/mem_reg[6][8]  ( .D(n2226), .CK(clk), .QN(\mx/mem[6][8] ) );
  DFF_X1 \mx/mem_reg[6][7]  ( .D(n2225), .CK(clk), .QN(\mx/mem[6][7] ) );
  DFF_X1 \mx/mem_reg[6][6]  ( .D(n2224), .CK(clk), .QN(\mx/mem[6][6] ) );
  DFF_X1 \mx/mem_reg[6][5]  ( .D(n2223), .CK(clk), .QN(\mx/mem[6][5] ) );
  DFF_X1 \mx/mem_reg[6][4]  ( .D(n2222), .CK(clk), .QN(\mx/mem[6][4] ) );
  DFF_X1 \mx/mem_reg[6][3]  ( .D(n2221), .CK(clk), .QN(\mx/mem[6][3] ) );
  DFF_X1 \mx/mem_reg[6][2]  ( .D(n2220), .CK(clk), .QN(\mx/mem[6][2] ) );
  DFF_X1 \mx/mem_reg[6][1]  ( .D(n2219), .CK(clk), .QN(\mx/mem[6][1] ) );
  DFF_X1 \mx/mem_reg[6][0]  ( .D(n2218), .CK(clk), .QN(\mx/mem[6][0] ) );
  DFF_X1 \mx/mem_reg[15][15]  ( .D(n2377), .CK(clk), .QN(\mx/mem[15][15] ) );
  DFF_X1 \mx/mem_reg[15][14]  ( .D(n2376), .CK(clk), .QN(\mx/mem[15][14] ) );
  DFF_X1 \mx/mem_reg[15][13]  ( .D(n2375), .CK(clk), .QN(\mx/mem[15][13] ) );
  DFF_X1 \mx/mem_reg[15][12]  ( .D(n2374), .CK(clk), .QN(\mx/mem[15][12] ) );
  DFF_X1 \mx/mem_reg[15][11]  ( .D(n2373), .CK(clk), .QN(\mx/mem[15][11] ) );
  DFF_X1 \mx/mem_reg[15][10]  ( .D(n2372), .CK(clk), .QN(\mx/mem[15][10] ) );
  DFF_X1 \mx/mem_reg[15][9]  ( .D(n2371), .CK(clk), .QN(\mx/mem[15][9] ) );
  DFF_X1 \mx/mem_reg[15][8]  ( .D(n2370), .CK(clk), .QN(\mx/mem[15][8] ) );
  DFF_X1 \mx/mem_reg[15][7]  ( .D(n2369), .CK(clk), .QN(\mx/mem[15][7] ) );
  DFF_X1 \mx/mem_reg[15][6]  ( .D(n2368), .CK(clk), .QN(\mx/mem[15][6] ) );
  DFF_X1 \mx/mem_reg[15][5]  ( .D(n2367), .CK(clk), .QN(\mx/mem[15][5] ) );
  DFF_X1 \mx/mem_reg[15][4]  ( .D(n2366), .CK(clk), .QN(\mx/mem[15][4] ) );
  DFF_X1 \mx/mem_reg[15][3]  ( .D(n2365), .CK(clk), .QN(\mx/mem[15][3] ) );
  DFF_X1 \mx/mem_reg[15][2]  ( .D(n2364), .CK(clk), .QN(\mx/mem[15][2] ) );
  DFF_X1 \mx/mem_reg[15][1]  ( .D(n2363), .CK(clk), .QN(\mx/mem[15][1] ) );
  DFF_X1 \mx/mem_reg[15][0]  ( .D(n2362), .CK(clk), .QN(\mx/mem[15][0] ) );
  DFF_X1 \mx/mem_reg[14][15]  ( .D(n2361), .CK(clk), .QN(\mx/mem[14][15] ) );
  DFF_X1 \mx/mem_reg[14][14]  ( .D(n2360), .CK(clk), .QN(\mx/mem[14][14] ) );
  DFF_X1 \mx/mem_reg[14][13]  ( .D(n2359), .CK(clk), .QN(\mx/mem[14][13] ) );
  DFF_X1 \mx/mem_reg[14][12]  ( .D(n2358), .CK(clk), .QN(\mx/mem[14][12] ) );
  DFF_X1 \mx/mem_reg[14][11]  ( .D(n2357), .CK(clk), .QN(\mx/mem[14][11] ) );
  DFF_X1 \mx/mem_reg[14][10]  ( .D(n2356), .CK(clk), .QN(\mx/mem[14][10] ) );
  DFF_X1 \mx/mem_reg[14][9]  ( .D(n2355), .CK(clk), .QN(\mx/mem[14][9] ) );
  DFF_X1 \mx/mem_reg[14][8]  ( .D(n2354), .CK(clk), .QN(\mx/mem[14][8] ) );
  DFF_X1 \mx/mem_reg[14][7]  ( .D(n2353), .CK(clk), .QN(\mx/mem[14][7] ) );
  DFF_X1 \mx/mem_reg[14][6]  ( .D(n2352), .CK(clk), .QN(\mx/mem[14][6] ) );
  DFF_X1 \mx/mem_reg[14][5]  ( .D(n2351), .CK(clk), .QN(\mx/mem[14][5] ) );
  DFF_X1 \mx/mem_reg[14][4]  ( .D(n2350), .CK(clk), .QN(\mx/mem[14][4] ) );
  DFF_X1 \mx/mem_reg[14][3]  ( .D(n2349), .CK(clk), .QN(\mx/mem[14][3] ) );
  DFF_X1 \mx/mem_reg[14][2]  ( .D(n2348), .CK(clk), .QN(\mx/mem[14][2] ) );
  DFF_X1 \mx/mem_reg[14][1]  ( .D(n2347), .CK(clk), .QN(\mx/mem[14][1] ) );
  DFF_X1 \mx/mem_reg[14][0]  ( .D(n2346), .CK(clk), .QN(\mx/mem[14][0] ) );
  DFF_X1 \mx/mem_reg[7][15]  ( .D(n2249), .CK(clk), .QN(\mx/mem[7][15] ) );
  DFF_X1 \mx/mem_reg[7][14]  ( .D(n2248), .CK(clk), .QN(\mx/mem[7][14] ) );
  DFF_X1 \mx/mem_reg[7][13]  ( .D(n2247), .CK(clk), .QN(\mx/mem[7][13] ) );
  DFF_X1 \mx/mem_reg[7][12]  ( .D(n2246), .CK(clk), .QN(\mx/mem[7][12] ) );
  DFF_X1 \mx/mem_reg[7][11]  ( .D(n2245), .CK(clk), .QN(\mx/mem[7][11] ) );
  DFF_X1 \mx/mem_reg[7][10]  ( .D(n2244), .CK(clk), .QN(\mx/mem[7][10] ) );
  DFF_X1 \mx/mem_reg[7][9]  ( .D(n2243), .CK(clk), .QN(\mx/mem[7][9] ) );
  DFF_X1 \mx/mem_reg[7][8]  ( .D(n2242), .CK(clk), .QN(\mx/mem[7][8] ) );
  DFF_X1 \mx/mem_reg[7][7]  ( .D(n2241), .CK(clk), .QN(\mx/mem[7][7] ) );
  DFF_X1 \mx/mem_reg[7][6]  ( .D(n2240), .CK(clk), .QN(\mx/mem[7][6] ) );
  DFF_X1 \mx/mem_reg[7][5]  ( .D(n2239), .CK(clk), .QN(\mx/mem[7][5] ) );
  DFF_X1 \mx/mem_reg[7][4]  ( .D(n2238), .CK(clk), .QN(\mx/mem[7][4] ) );
  DFF_X1 \mx/mem_reg[7][3]  ( .D(n2237), .CK(clk), .QN(\mx/mem[7][3] ) );
  DFF_X1 \mx/mem_reg[7][2]  ( .D(n2236), .CK(clk), .QN(\mx/mem[7][2] ) );
  DFF_X1 \mx/mem_reg[7][1]  ( .D(n2235), .CK(clk), .QN(\mx/mem[7][1] ) );
  DFF_X1 \mx/mem_reg[7][0]  ( .D(n2234), .CK(clk), .QN(\mx/mem[7][0] ) );
  DFF_X1 \mx/mem_reg[9][15]  ( .D(n2281), .CK(clk), .QN(\mx/mem[9][15] ) );
  DFF_X1 \mx/mem_reg[9][14]  ( .D(n2280), .CK(clk), .QN(\mx/mem[9][14] ) );
  DFF_X1 \mx/mem_reg[9][13]  ( .D(n2279), .CK(clk), .QN(\mx/mem[9][13] ) );
  DFF_X1 \mx/mem_reg[9][12]  ( .D(n2278), .CK(clk), .QN(\mx/mem[9][12] ) );
  DFF_X1 \mx/mem_reg[9][11]  ( .D(n2277), .CK(clk), .QN(\mx/mem[9][11] ) );
  DFF_X1 \mx/mem_reg[9][10]  ( .D(n2276), .CK(clk), .QN(\mx/mem[9][10] ) );
  DFF_X1 \mx/mem_reg[9][9]  ( .D(n2275), .CK(clk), .QN(\mx/mem[9][9] ) );
  DFF_X1 \mx/mem_reg[9][8]  ( .D(n2274), .CK(clk), .QN(\mx/mem[9][8] ) );
  DFF_X1 \mx/mem_reg[9][7]  ( .D(n2273), .CK(clk), .QN(\mx/mem[9][7] ) );
  DFF_X1 \mx/mem_reg[9][6]  ( .D(n2272), .CK(clk), .QN(\mx/mem[9][6] ) );
  DFF_X1 \mx/mem_reg[9][5]  ( .D(n2271), .CK(clk), .QN(\mx/mem[9][5] ) );
  DFF_X1 \mx/mem_reg[9][4]  ( .D(n2270), .CK(clk), .QN(\mx/mem[9][4] ) );
  DFF_X1 \mx/mem_reg[9][3]  ( .D(n2269), .CK(clk), .QN(\mx/mem[9][3] ) );
  DFF_X1 \mx/mem_reg[9][2]  ( .D(n2268), .CK(clk), .QN(\mx/mem[9][2] ) );
  DFF_X1 \mx/mem_reg[9][1]  ( .D(n2267), .CK(clk), .QN(\mx/mem[9][1] ) );
  DFF_X1 \mx/mem_reg[9][0]  ( .D(n2266), .CK(clk), .QN(\mx/mem[9][0] ) );
  DFF_X1 \mx/mem_reg[8][15]  ( .D(n2265), .CK(clk), .QN(\mx/mem[8][15] ) );
  DFF_X1 \mx/mem_reg[8][14]  ( .D(n2264), .CK(clk), .QN(\mx/mem[8][14] ) );
  DFF_X1 \mx/mem_reg[8][13]  ( .D(n2263), .CK(clk), .QN(\mx/mem[8][13] ) );
  DFF_X1 \mx/mem_reg[8][12]  ( .D(n2262), .CK(clk), .QN(\mx/mem[8][12] ) );
  DFF_X1 \mx/mem_reg[8][11]  ( .D(n2261), .CK(clk), .QN(\mx/mem[8][11] ) );
  DFF_X1 \mx/mem_reg[8][10]  ( .D(n2260), .CK(clk), .QN(\mx/mem[8][10] ) );
  DFF_X1 \mx/mem_reg[8][9]  ( .D(n2259), .CK(clk), .QN(\mx/mem[8][9] ) );
  DFF_X1 \mx/mem_reg[8][8]  ( .D(n2258), .CK(clk), .QN(\mx/mem[8][8] ) );
  DFF_X1 \mx/mem_reg[8][7]  ( .D(n2257), .CK(clk), .QN(\mx/mem[8][7] ) );
  DFF_X1 \mx/mem_reg[8][6]  ( .D(n2256), .CK(clk), .QN(\mx/mem[8][6] ) );
  DFF_X1 \mx/mem_reg[8][5]  ( .D(n2255), .CK(clk), .QN(\mx/mem[8][5] ) );
  DFF_X1 \mx/mem_reg[8][4]  ( .D(n2254), .CK(clk), .QN(\mx/mem[8][4] ) );
  DFF_X1 \mx/mem_reg[8][3]  ( .D(n2253), .CK(clk), .QN(\mx/mem[8][3] ) );
  DFF_X1 \mx/mem_reg[8][2]  ( .D(n2252), .CK(clk), .QN(\mx/mem[8][2] ) );
  DFF_X1 \mx/mem_reg[8][1]  ( .D(n2251), .CK(clk), .QN(\mx/mem[8][1] ) );
  DFF_X1 \mx/mem_reg[8][0]  ( .D(n2250), .CK(clk), .QN(\mx/mem[8][0] ) );
  DFF_X1 \mx/mem_reg[1][15]  ( .D(n2153), .CK(clk), .QN(\mx/mem[1][15] ) );
  DFF_X1 \mx/mem_reg[1][14]  ( .D(n2152), .CK(clk), .QN(\mx/mem[1][14] ) );
  DFF_X1 \mx/mem_reg[1][13]  ( .D(n2151), .CK(clk), .QN(\mx/mem[1][13] ) );
  DFF_X1 \mx/mem_reg[1][12]  ( .D(n2150), .CK(clk), .QN(\mx/mem[1][12] ) );
  DFF_X1 \mx/mem_reg[1][11]  ( .D(n2149), .CK(clk), .QN(\mx/mem[1][11] ) );
  DFF_X1 \mx/mem_reg[1][10]  ( .D(n2148), .CK(clk), .QN(\mx/mem[1][10] ) );
  DFF_X1 \mx/mem_reg[1][9]  ( .D(n2147), .CK(clk), .QN(\mx/mem[1][9] ) );
  DFF_X1 \mx/mem_reg[1][8]  ( .D(n2146), .CK(clk), .QN(\mx/mem[1][8] ) );
  DFF_X1 \mx/mem_reg[1][7]  ( .D(n2145), .CK(clk), .QN(\mx/mem[1][7] ) );
  DFF_X1 \mx/mem_reg[1][6]  ( .D(n2144), .CK(clk), .QN(\mx/mem[1][6] ) );
  DFF_X1 \mx/mem_reg[1][5]  ( .D(n2143), .CK(clk), .QN(\mx/mem[1][5] ) );
  DFF_X1 \mx/mem_reg[1][4]  ( .D(n2142), .CK(clk), .QN(\mx/mem[1][4] ) );
  DFF_X1 \mx/mem_reg[1][3]  ( .D(n2141), .CK(clk), .QN(\mx/mem[1][3] ) );
  DFF_X1 \mx/mem_reg[1][2]  ( .D(n2140), .CK(clk), .QN(\mx/mem[1][2] ) );
  DFF_X1 \mx/mem_reg[1][1]  ( .D(n2139), .CK(clk), .QN(\mx/mem[1][1] ) );
  DFF_X1 \mx/mem_reg[1][0]  ( .D(n2138), .CK(clk), .QN(\mx/mem[1][0] ) );
  DFF_X1 \mx/mem_reg[0][15]  ( .D(n2137), .CK(clk), .QN(\mx/mem[0][15] ) );
  DFF_X1 \mx/mem_reg[0][14]  ( .D(n2136), .CK(clk), .QN(\mx/mem[0][14] ) );
  DFF_X1 \mx/mem_reg[0][13]  ( .D(n2135), .CK(clk), .QN(\mx/mem[0][13] ) );
  DFF_X1 \mx/mem_reg[0][12]  ( .D(n2134), .CK(clk), .QN(\mx/mem[0][12] ) );
  DFF_X1 \mx/mem_reg[0][11]  ( .D(n2133), .CK(clk), .QN(\mx/mem[0][11] ) );
  DFF_X1 \mx/mem_reg[0][10]  ( .D(n2132), .CK(clk), .QN(\mx/mem[0][10] ) );
  DFF_X1 \mx/mem_reg[0][9]  ( .D(n2131), .CK(clk), .QN(\mx/mem[0][9] ) );
  DFF_X1 \mx/mem_reg[0][8]  ( .D(n2130), .CK(clk), .QN(\mx/mem[0][8] ) );
  DFF_X1 \mx/mem_reg[0][7]  ( .D(n2129), .CK(clk), .QN(\mx/mem[0][7] ) );
  DFF_X1 \mx/mem_reg[0][6]  ( .D(n2128), .CK(clk), .QN(\mx/mem[0][6] ) );
  DFF_X1 \mx/mem_reg[0][5]  ( .D(n2127), .CK(clk), .QN(\mx/mem[0][5] ) );
  DFF_X1 \mx/mem_reg[0][4]  ( .D(n2126), .CK(clk), .QN(\mx/mem[0][4] ) );
  DFF_X1 \mx/mem_reg[0][3]  ( .D(n2125), .CK(clk), .QN(\mx/mem[0][3] ) );
  DFF_X1 \mx/mem_reg[0][2]  ( .D(n2124), .CK(clk), .QN(\mx/mem[0][2] ) );
  DFF_X1 \mx/mem_reg[0][1]  ( .D(n2123), .CK(clk), .QN(\mx/mem[0][1] ) );
  DFF_X1 \mx/mem_reg[0][0]  ( .D(n2122), .CK(clk), .QN(\mx/mem[0][0] ) );
  DFF_X1 \mx/mem_reg[11][15]  ( .D(n2313), .CK(clk), .QN(\mx/mem[11][15] ) );
  DFF_X1 \mx/mem_reg[11][14]  ( .D(n2312), .CK(clk), .QN(\mx/mem[11][14] ) );
  DFF_X1 \mx/mem_reg[11][13]  ( .D(n2311), .CK(clk), .QN(\mx/mem[11][13] ) );
  DFF_X1 \mx/mem_reg[11][12]  ( .D(n2310), .CK(clk), .QN(\mx/mem[11][12] ) );
  DFF_X1 \mx/mem_reg[11][11]  ( .D(n2309), .CK(clk), .QN(\mx/mem[11][11] ) );
  DFF_X1 \mx/mem_reg[11][10]  ( .D(n2308), .CK(clk), .QN(\mx/mem[11][10] ) );
  DFF_X1 \mx/mem_reg[11][9]  ( .D(n2307), .CK(clk), .QN(\mx/mem[11][9] ) );
  DFF_X1 \mx/mem_reg[11][8]  ( .D(n2306), .CK(clk), .QN(\mx/mem[11][8] ) );
  DFF_X1 \mx/mem_reg[11][7]  ( .D(n2305), .CK(clk), .QN(\mx/mem[11][7] ) );
  DFF_X1 \mx/mem_reg[11][6]  ( .D(n2304), .CK(clk), .QN(\mx/mem[11][6] ) );
  DFF_X1 \mx/mem_reg[11][5]  ( .D(n2303), .CK(clk), .QN(\mx/mem[11][5] ) );
  DFF_X1 \mx/mem_reg[11][4]  ( .D(n2302), .CK(clk), .QN(\mx/mem[11][4] ) );
  DFF_X1 \mx/mem_reg[11][3]  ( .D(n2301), .CK(clk), .QN(\mx/mem[11][3] ) );
  DFF_X1 \mx/mem_reg[11][2]  ( .D(n2300), .CK(clk), .QN(\mx/mem[11][2] ) );
  DFF_X1 \mx/mem_reg[11][1]  ( .D(n2299), .CK(clk), .QN(\mx/mem[11][1] ) );
  DFF_X1 \mx/mem_reg[11][0]  ( .D(n2298), .CK(clk), .QN(\mx/mem[11][0] ) );
  DFF_X1 \mx/mem_reg[10][15]  ( .D(n2297), .CK(clk), .QN(\mx/mem[10][15] ) );
  DFF_X1 \mx/mem_reg[10][14]  ( .D(n2296), .CK(clk), .QN(\mx/mem[10][14] ) );
  DFF_X1 \mx/mem_reg[10][13]  ( .D(n2295), .CK(clk), .QN(\mx/mem[10][13] ) );
  DFF_X1 \mx/mem_reg[10][12]  ( .D(n2294), .CK(clk), .QN(\mx/mem[10][12] ) );
  DFF_X1 \mx/mem_reg[10][11]  ( .D(n2293), .CK(clk), .QN(\mx/mem[10][11] ) );
  DFF_X1 \mx/mem_reg[10][10]  ( .D(n2292), .CK(clk), .QN(\mx/mem[10][10] ) );
  DFF_X1 \mx/mem_reg[10][9]  ( .D(n2291), .CK(clk), .QN(\mx/mem[10][9] ) );
  DFF_X1 \mx/mem_reg[10][8]  ( .D(n2290), .CK(clk), .QN(\mx/mem[10][8] ) );
  DFF_X1 \mx/mem_reg[10][7]  ( .D(n2289), .CK(clk), .QN(\mx/mem[10][7] ) );
  DFF_X1 \mx/mem_reg[10][6]  ( .D(n2288), .CK(clk), .QN(\mx/mem[10][6] ) );
  DFF_X1 \mx/mem_reg[10][5]  ( .D(n2287), .CK(clk), .QN(\mx/mem[10][5] ) );
  DFF_X1 \mx/mem_reg[10][4]  ( .D(n2286), .CK(clk), .QN(\mx/mem[10][4] ) );
  DFF_X1 \mx/mem_reg[10][3]  ( .D(n2285), .CK(clk), .QN(\mx/mem[10][3] ) );
  DFF_X1 \mx/mem_reg[10][2]  ( .D(n2284), .CK(clk), .QN(\mx/mem[10][2] ) );
  DFF_X1 \mx/mem_reg[10][1]  ( .D(n2283), .CK(clk), .QN(\mx/mem[10][1] ) );
  DFF_X1 \mx/mem_reg[10][0]  ( .D(n2282), .CK(clk), .QN(\mx/mem[10][0] ) );
  DFF_X1 \mx/mem_reg[3][15]  ( .D(n2185), .CK(clk), .QN(\mx/mem[3][15] ) );
  DFF_X1 \mx/mem_reg[3][14]  ( .D(n2184), .CK(clk), .QN(\mx/mem[3][14] ) );
  DFF_X1 \mx/mem_reg[3][13]  ( .D(n2183), .CK(clk), .QN(\mx/mem[3][13] ) );
  DFF_X1 \mx/mem_reg[3][12]  ( .D(n2182), .CK(clk), .QN(\mx/mem[3][12] ) );
  DFF_X1 \mx/mem_reg[3][11]  ( .D(n2181), .CK(clk), .QN(\mx/mem[3][11] ) );
  DFF_X1 \mx/mem_reg[3][10]  ( .D(n2180), .CK(clk), .QN(\mx/mem[3][10] ) );
  DFF_X1 \mx/mem_reg[3][9]  ( .D(n2179), .CK(clk), .QN(\mx/mem[3][9] ) );
  DFF_X1 \mx/mem_reg[3][8]  ( .D(n2178), .CK(clk), .QN(\mx/mem[3][8] ) );
  DFF_X1 \mx/mem_reg[3][7]  ( .D(n2177), .CK(clk), .QN(\mx/mem[3][7] ) );
  DFF_X1 \mx/mem_reg[3][6]  ( .D(n2176), .CK(clk), .QN(\mx/mem[3][6] ) );
  DFF_X1 \mx/mem_reg[3][5]  ( .D(n2175), .CK(clk), .QN(\mx/mem[3][5] ) );
  DFF_X1 \mx/mem_reg[3][4]  ( .D(n2174), .CK(clk), .QN(\mx/mem[3][4] ) );
  DFF_X1 \mx/mem_reg[3][3]  ( .D(n2173), .CK(clk), .QN(\mx/mem[3][3] ) );
  DFF_X1 \mx/mem_reg[3][2]  ( .D(n2172), .CK(clk), .QN(\mx/mem[3][2] ) );
  DFF_X1 \mx/mem_reg[3][1]  ( .D(n2171), .CK(clk), .QN(\mx/mem[3][1] ) );
  DFF_X1 \mx/mem_reg[3][0]  ( .D(n2170), .CK(clk), .QN(\mx/mem[3][0] ) );
  DFF_X1 \mx/mem_reg[2][15]  ( .D(n2169), .CK(clk), .QN(\mx/mem[2][15] ) );
  DFF_X1 \mx/mem_reg[2][14]  ( .D(n2168), .CK(clk), .QN(\mx/mem[2][14] ) );
  DFF_X1 \mx/mem_reg[2][13]  ( .D(n2167), .CK(clk), .QN(\mx/mem[2][13] ) );
  DFF_X1 \mx/mem_reg[2][12]  ( .D(n2166), .CK(clk), .QN(\mx/mem[2][12] ) );
  DFF_X1 \mx/mem_reg[2][11]  ( .D(n2165), .CK(clk), .QN(\mx/mem[2][11] ) );
  DFF_X1 \mx/mem_reg[2][10]  ( .D(n2164), .CK(clk), .QN(\mx/mem[2][10] ) );
  DFF_X1 \mx/mem_reg[2][9]  ( .D(n2163), .CK(clk), .QN(\mx/mem[2][9] ) );
  DFF_X1 \mx/mem_reg[2][8]  ( .D(n2162), .CK(clk), .QN(\mx/mem[2][8] ) );
  DFF_X1 \mx/mem_reg[2][7]  ( .D(n2161), .CK(clk), .QN(\mx/mem[2][7] ) );
  DFF_X1 \mx/mem_reg[2][6]  ( .D(n2160), .CK(clk), .QN(\mx/mem[2][6] ) );
  DFF_X1 \mx/mem_reg[2][5]  ( .D(n2159), .CK(clk), .QN(\mx/mem[2][5] ) );
  DFF_X1 \mx/mem_reg[2][4]  ( .D(n2158), .CK(clk), .QN(\mx/mem[2][4] ) );
  DFF_X1 \mx/mem_reg[2][3]  ( .D(n2157), .CK(clk), .QN(\mx/mem[2][3] ) );
  DFF_X1 \mx/mem_reg[2][2]  ( .D(n2156), .CK(clk), .QN(\mx/mem[2][2] ) );
  DFF_X1 \mx/mem_reg[2][1]  ( .D(n2155), .CK(clk), .QN(\mx/mem[2][1] ) );
  DFF_X1 \mx/mem_reg[2][0]  ( .D(n2154), .CK(clk), .QN(\mx/mem[2][0] ) );
  DFF_X1 \mx/mem_reg[13][15]  ( .D(n2345), .CK(clk), .QN(\mx/mem[13][15] ) );
  DFF_X1 \mx/mem_reg[13][14]  ( .D(n2344), .CK(clk), .QN(\mx/mem[13][14] ) );
  DFF_X1 \mx/mem_reg[13][13]  ( .D(n2343), .CK(clk), .QN(\mx/mem[13][13] ) );
  DFF_X1 \mx/mem_reg[13][12]  ( .D(n2342), .CK(clk), .QN(\mx/mem[13][12] ) );
  DFF_X1 \mx/mem_reg[13][11]  ( .D(n2341), .CK(clk), .QN(\mx/mem[13][11] ) );
  DFF_X1 \mx/mem_reg[13][10]  ( .D(n2340), .CK(clk), .QN(\mx/mem[13][10] ) );
  DFF_X1 \mx/mem_reg[13][9]  ( .D(n2339), .CK(clk), .QN(\mx/mem[13][9] ) );
  DFF_X1 \mx/mem_reg[13][8]  ( .D(n2338), .CK(clk), .QN(\mx/mem[13][8] ) );
  DFF_X1 \mx/mem_reg[13][7]  ( .D(n2337), .CK(clk), .QN(\mx/mem[13][7] ) );
  DFF_X1 \mx/mem_reg[13][6]  ( .D(n2336), .CK(clk), .QN(\mx/mem[13][6] ) );
  DFF_X1 \mx/mem_reg[13][5]  ( .D(n2335), .CK(clk), .QN(\mx/mem[13][5] ) );
  DFF_X1 \mx/mem_reg[13][4]  ( .D(n2334), .CK(clk), .QN(\mx/mem[13][4] ) );
  DFF_X1 \mx/mem_reg[13][3]  ( .D(n2333), .CK(clk), .QN(\mx/mem[13][3] ) );
  DFF_X1 \mx/mem_reg[13][2]  ( .D(n2332), .CK(clk), .QN(\mx/mem[13][2] ) );
  DFF_X1 \mx/mem_reg[13][1]  ( .D(n2331), .CK(clk), .QN(\mx/mem[13][1] ) );
  DFF_X1 \mx/mem_reg[13][0]  ( .D(n2330), .CK(clk), .QN(\mx/mem[13][0] ) );
  DFF_X1 \mx/mem_reg[12][15]  ( .D(n2329), .CK(clk), .QN(\mx/mem[12][15] ) );
  DFF_X1 \mx/mem_reg[12][14]  ( .D(n2328), .CK(clk), .QN(\mx/mem[12][14] ) );
  DFF_X1 \mx/mem_reg[12][13]  ( .D(n2327), .CK(clk), .QN(\mx/mem[12][13] ) );
  DFF_X1 \mx/mem_reg[12][12]  ( .D(n2326), .CK(clk), .QN(\mx/mem[12][12] ) );
  DFF_X1 \mx/mem_reg[12][11]  ( .D(n2325), .CK(clk), .QN(\mx/mem[12][11] ) );
  DFF_X1 \mx/mem_reg[12][10]  ( .D(n2324), .CK(clk), .QN(\mx/mem[12][10] ) );
  DFF_X1 \mx/mem_reg[12][9]  ( .D(n2323), .CK(clk), .QN(\mx/mem[12][9] ) );
  DFF_X1 \mx/mem_reg[12][8]  ( .D(n2322), .CK(clk), .QN(\mx/mem[12][8] ) );
  DFF_X1 \mx/mem_reg[12][7]  ( .D(n2321), .CK(clk), .QN(\mx/mem[12][7] ) );
  DFF_X1 \mx/mem_reg[12][6]  ( .D(n2320), .CK(clk), .QN(\mx/mem[12][6] ) );
  DFF_X1 \mx/mem_reg[12][5]  ( .D(n2319), .CK(clk), .QN(\mx/mem[12][5] ) );
  DFF_X1 \mx/mem_reg[12][4]  ( .D(n2318), .CK(clk), .QN(\mx/mem[12][4] ) );
  DFF_X1 \mx/mem_reg[12][3]  ( .D(n2317), .CK(clk), .QN(\mx/mem[12][3] ) );
  DFF_X1 \mx/mem_reg[12][2]  ( .D(n2316), .CK(clk), .QN(\mx/mem[12][2] ) );
  DFF_X1 \mx/mem_reg[12][1]  ( .D(n2315), .CK(clk), .QN(\mx/mem[12][1] ) );
  DFF_X1 \mx/mem_reg[12][0]  ( .D(n2314), .CK(clk), .QN(\mx/mem[12][0] ) );
  DFF_X1 \mx/mem_reg[5][15]  ( .D(n2217), .CK(clk), .QN(\mx/mem[5][15] ) );
  DFF_X1 \mx/mem_reg[5][14]  ( .D(n2216), .CK(clk), .QN(\mx/mem[5][14] ) );
  DFF_X1 \mx/mem_reg[5][13]  ( .D(n2215), .CK(clk), .QN(\mx/mem[5][13] ) );
  DFF_X1 \mx/mem_reg[5][12]  ( .D(n2214), .CK(clk), .QN(\mx/mem[5][12] ) );
  DFF_X1 \mx/mem_reg[5][11]  ( .D(n2213), .CK(clk), .QN(\mx/mem[5][11] ) );
  DFF_X1 \mx/mem_reg[5][10]  ( .D(n2212), .CK(clk), .QN(\mx/mem[5][10] ) );
  DFF_X1 \mx/mem_reg[5][9]  ( .D(n2211), .CK(clk), .QN(\mx/mem[5][9] ) );
  DFF_X1 \mx/mem_reg[5][8]  ( .D(n2210), .CK(clk), .QN(\mx/mem[5][8] ) );
  DFF_X1 \mx/mem_reg[5][7]  ( .D(n2209), .CK(clk), .QN(\mx/mem[5][7] ) );
  DFF_X1 \mx/mem_reg[5][6]  ( .D(n2208), .CK(clk), .QN(\mx/mem[5][6] ) );
  DFF_X1 \mx/mem_reg[5][5]  ( .D(n2207), .CK(clk), .QN(\mx/mem[5][5] ) );
  DFF_X1 \mx/mem_reg[5][4]  ( .D(n2206), .CK(clk), .QN(\mx/mem[5][4] ) );
  DFF_X1 \mx/mem_reg[5][3]  ( .D(n2205), .CK(clk), .QN(\mx/mem[5][3] ) );
  DFF_X1 \mx/mem_reg[5][2]  ( .D(n2204), .CK(clk), .QN(\mx/mem[5][2] ) );
  DFF_X1 \mx/mem_reg[5][1]  ( .D(n2203), .CK(clk), .QN(\mx/mem[5][1] ) );
  DFF_X1 \mx/mem_reg[5][0]  ( .D(n2202), .CK(clk), .QN(\mx/mem[5][0] ) );
  DFF_X1 \mx/mem_reg[4][15]  ( .D(n2201), .CK(clk), .QN(\mx/mem[4][15] ) );
  DFF_X1 \mx/mem_reg[4][14]  ( .D(n2200), .CK(clk), .QN(\mx/mem[4][14] ) );
  DFF_X1 \mx/mem_reg[4][13]  ( .D(n2199), .CK(clk), .QN(\mx/mem[4][13] ) );
  DFF_X1 \mx/mem_reg[4][12]  ( .D(n2198), .CK(clk), .QN(\mx/mem[4][12] ) );
  DFF_X1 \mx/mem_reg[4][11]  ( .D(n2197), .CK(clk), .QN(\mx/mem[4][11] ) );
  DFF_X1 \mx/mem_reg[4][10]  ( .D(n2196), .CK(clk), .QN(\mx/mem[4][10] ) );
  DFF_X1 \mx/mem_reg[4][9]  ( .D(n2195), .CK(clk), .QN(\mx/mem[4][9] ) );
  DFF_X1 \mx/mem_reg[4][8]  ( .D(n2194), .CK(clk), .QN(\mx/mem[4][8] ) );
  DFF_X1 \mx/mem_reg[4][7]  ( .D(n2193), .CK(clk), .QN(\mx/mem[4][7] ) );
  DFF_X1 \mx/mem_reg[4][6]  ( .D(n2192), .CK(clk), .QN(\mx/mem[4][6] ) );
  DFF_X1 \mx/mem_reg[4][5]  ( .D(n2191), .CK(clk), .QN(\mx/mem[4][5] ) );
  DFF_X1 \mx/mem_reg[4][4]  ( .D(n2190), .CK(clk), .QN(\mx/mem[4][4] ) );
  DFF_X1 \mx/mem_reg[4][3]  ( .D(n2189), .CK(clk), .QN(\mx/mem[4][3] ) );
  DFF_X1 \mx/mem_reg[4][2]  ( .D(n2188), .CK(clk), .QN(\mx/mem[4][2] ) );
  DFF_X1 \mx/mem_reg[4][1]  ( .D(n2187), .CK(clk), .QN(\mx/mem[4][1] ) );
  DFF_X1 \mx/mem_reg[4][0]  ( .D(n2186), .CK(clk), .QN(\mx/mem[4][0] ) );
  DFF_X1 \mx/data_out_reg[2]  ( .D(n1012), .CK(clk), .QN(w_to_multx[2]) );
  DFF_X1 \conv/prev_output_reg[15]  ( .D(\conv/N125 ), .CK(clk), .QN(n2099) );
  DFFRS_X1 \conv/prev_output_reg[3]  ( .D(\conv/N113 ), .CK(clk), .RN(1'b1), 
        .SN(1'b1), .Q(n2101) );
  DFF_X1 \mx/data_out_reg[11]  ( .D(\mx/N18 ), .CK(clk), .Q(n964), .QN(n1016)
         );
  DFF_X2 \mf/z_reg[1]  ( .D(\mf/N12 ), .CK(clk), .Q(w_to_multf[1]), .QN(n962)
         );
  DFF_X1 \conv/m_data_out_y_reg[14]  ( .D(\conv/N146 ), .CK(clk), .Q(
        m_data_out_y[14]) );
  DFF_X1 \mx/data_out_reg[13]  ( .D(\mx/N16 ), .CK(clk), .Q(w_to_multx[13]), 
        .QN(n1015) );
  DFF_X1 \mx/data_out_reg[3]  ( .D(\mx/N26 ), .CK(clk), .Q(w_to_multx[3]), 
        .QN(n1017) );
  DFF_X1 \conv/m_data_out_y_reg[8]  ( .D(\conv/N140 ), .CK(clk), .Q(
        m_data_out_y[8]) );
  DFF_X1 \conv/m_data_out_y_reg[5]  ( .D(\conv/N137 ), .CK(clk), .Q(
        m_data_out_y[5]) );
  DFF_X1 \conv/m_data_out_y_reg[10]  ( .D(\conv/N142 ), .CK(clk), .Q(
        m_data_out_y[10]) );
  DFF_X1 \conv/m_data_out_y_reg[11]  ( .D(\conv/N143 ), .CK(clk), .Q(
        m_data_out_y[11]) );
  DFF_X1 \conv/m_data_out_y_reg[3]  ( .D(\conv/N135 ), .CK(clk), .Q(
        m_data_out_y[3]) );
  DFF_X1 \conv/m_data_out_y_reg[12]  ( .D(\conv/N144 ), .CK(clk), .Q(
        m_data_out_y[12]) );
  DFF_X1 \conv/m_data_out_y_reg[1]  ( .D(\conv/N133 ), .CK(clk), .Q(
        m_data_out_y[1]) );
  DFF_X1 \conv/m_data_out_y_reg[2]  ( .D(\conv/N134 ), .CK(clk), .Q(
        m_data_out_y[2]) );
  DFF_X1 \conv/m_data_out_y_reg[0]  ( .D(\conv/N132 ), .CK(clk), .Q(
        m_data_out_y[0]) );
  DFF_X1 \conv/m_data_out_y_reg[6]  ( .D(\conv/N138 ), .CK(clk), .Q(
        m_data_out_y[6]) );
  DFF_X1 \conv/m_data_out_y_reg[4]  ( .D(\conv/N136 ), .CK(clk), .Q(
        m_data_out_y[4]) );
  DFF_X1 \mf/z_reg[4]  ( .D(\mf/N14 ), .CK(clk), .Q(w_to_multf[4]), .QN(n968)
         );
  DFF_X1 \mf/z_reg[2]  ( .D(\mf/N13 ), .CK(clk), .Q(w_to_multf[2]), .QN(n959)
         );
  DFF_X1 \conv/prev_output_reg[8]  ( .D(\conv/N118 ), .CK(clk), .Q(
        \conv/prev_output [8]) );
  DFF_X1 \conv/prev_output_reg[7]  ( .D(\conv/N117 ), .CK(clk), .Q(
        \conv/prev_output [7]) );
  DFF_X1 \conv/prev_output_reg[6]  ( .D(\conv/N116 ), .CK(clk), .Q(
        \conv/prev_output [6]) );
  DFF_X1 \conv/prev_output_reg[5]  ( .D(\conv/N115 ), .CK(clk), .Q(
        \conv/prev_output [5]), .QN(n2102) );
  DFF_X1 \conv/prev_output_reg[4]  ( .D(\conv/N114 ), .CK(clk), .Q(
        \conv/prev_output [4]) );
  DFF_X1 \conv/prev_output_reg[2]  ( .D(\conv/N112 ), .CK(clk), .Q(
        \conv/prev_output [2]) );
  DFF_X1 \conv/prev_output_reg[1]  ( .D(\conv/N111 ), .CK(clk), .Q(
        \conv/prev_output [1]) );
  DFF_X1 \conv/prev_output_reg[0]  ( .D(\conv/N110 ), .CK(clk), .Q(
        \conv/prev_output [0]) );
  DFF_X1 \conv/prev_output_reg[14]  ( .D(\conv/N124 ), .CK(clk), .Q(
        \conv/prev_output [14]), .QN(n2098) );
  DFF_X1 \conv/prev_output_reg[9]  ( .D(\conv/N119 ), .CK(clk), .Q(
        \conv/prev_output [9]), .QN(n2103) );
  DFF_X1 \conv/prev_output_reg[12]  ( .D(\conv/N122 ), .CK(clk), .Q(
        \conv/prev_output [12]) );
  DFF_X1 \conv/prev_output_reg[13]  ( .D(\conv/N123 ), .CK(clk), .Q(
        \conv/prev_output [13]) );
  DFF_X1 \conv/prev_output_reg[10]  ( .D(\conv/N120 ), .CK(clk), .Q(
        \conv/prev_output [10]) );
  DFF_X1 \mx/data_out_reg[0]  ( .D(\mx/N29 ), .CK(clk), .Q(w_to_multx[0]), 
        .QN(n2105) );
  AOI21_X1 U1002 ( .B1(n1337), .B2(n1336), .A(n1335), .ZN(n1338) );
  NAND2_X1 U1003 ( .A1(n933), .A2(n932), .ZN(n1332) );
  OAI21_X1 U1004 ( .B1(n1305), .B2(n1304), .A(n934), .ZN(n933) );
  NAND2_X1 U1005 ( .A1(n931), .A2(n930), .ZN(n1325) );
  OAI21_X1 U1006 ( .B1(n1298), .B2(n1299), .A(n1297), .ZN(n931) );
  BUF_X1 U1007 ( .A(n1131), .Z(n1259) );
  NAND2_X1 U1008 ( .A1(n1101), .A2(n965), .ZN(n971) );
  XNOR2_X1 U1009 ( .A(n2104), .B(n968), .ZN(n1271) );
  NAND2_X2 U1010 ( .A1(n1299), .A2(n1298), .ZN(n930) );
  NAND2_X2 U1011 ( .A1(n1305), .A2(n1304), .ZN(n932) );
  XNOR2_X1 U1012 ( .A(n936), .B(n934), .ZN(n1608) );
  XNOR2_X1 U1013 ( .A(n935), .B(n1297), .ZN(n934) );
  XNOR2_X1 U1014 ( .A(n1299), .B(n1298), .ZN(n935) );
  XNOR2_X1 U1015 ( .A(n1305), .B(n1304), .ZN(n936) );
  AND2_X2 U1016 ( .A1(n1803), .A2(n1802), .ZN(n1005) );
  XNOR2_X1 U1017 ( .A(n937), .B(n1022), .ZN(n1101) );
  INV_X1 U1018 ( .A(n1016), .ZN(n937) );
  OAI21_X1 U1019 ( .B1(n1881), .B2(n1884), .A(n1885), .ZN(n1653) );
  NAND2_X1 U1020 ( .A1(n1639), .A2(\conv/prev_output [8]), .ZN(n1881) );
  NAND2_X1 U1021 ( .A1(n938), .A2(n1344), .ZN(n1385) );
  NAND2_X1 U1022 ( .A1(n1342), .A2(n1341), .ZN(n938) );
  BUF_X2 U1023 ( .A(n1131), .Z(n1276) );
  BUF_X1 U1024 ( .A(n1100), .Z(n1404) );
  OR2_X1 U1025 ( .A1(n1601), .A2(n1600), .ZN(n1603) );
  NAND2_X1 U1026 ( .A1(n1189), .A2(n1188), .ZN(n1585) );
  AND2_X2 U1027 ( .A1(n989), .A2(n1525), .ZN(n988) );
  BUF_X2 U1028 ( .A(n1094), .Z(n1400) );
  AND3_X2 U1029 ( .A1(n1557), .A2(n1647), .A3(n2102), .ZN(n1785) );
  BUF_X2 U1030 ( .A(n1100), .Z(n955) );
  BUF_X1 U1031 ( .A(n1584), .Z(n943) );
  BUF_X1 U1032 ( .A(w_to_multx[5]), .Z(n1213) );
  CLKBUF_X2 U1033 ( .A(w_to_multx[9]), .Z(n994) );
  CLKBUF_X2 U1034 ( .A(w_to_multf[7]), .Z(n951) );
  AND3_X1 U1035 ( .A1(n2111), .A2(e_acc), .A3(n1921), .ZN(n1804) );
  XNOR2_X1 U1036 ( .A(n1015), .B(n992), .ZN(n1505) );
  AND3_X1 U1037 ( .A1(n988), .A2(n1589), .A3(n2103), .ZN(n1884) );
  OR2_X1 U1038 ( .A1(n1241), .A2(n1240), .ZN(n1599) );
  AND2_X1 U1039 ( .A1(n1474), .A2(n1473), .ZN(n990) );
  OR2_X1 U1040 ( .A1(n1333), .A2(n1332), .ZN(n978) );
  OR2_X1 U1041 ( .A1(n1239), .A2(n1238), .ZN(n1569) );
  OR2_X1 U1042 ( .A1(n1180), .A2(n1179), .ZN(n1549) );
  AND2_X1 U1043 ( .A1(n1099), .A2(n1098), .ZN(n1422) );
  NAND2_X1 U1044 ( .A1(n1093), .A2(n1094), .ZN(n1402) );
  NAND2_X1 U1045 ( .A1(n1096), .A2(n1505), .ZN(n1504) );
  INV_X1 U1046 ( .A(n1039), .ZN(n973) );
  CLKBUF_X1 U1047 ( .A(n964), .Z(n945) );
  INV_X1 U1048 ( .A(n1017), .ZN(n979) );
  INV_X1 U1049 ( .A(n1505), .ZN(n939) );
  CLKBUF_X1 U1050 ( .A(n2378), .Z(n969) );
  NOR2_X1 U1051 ( .A1(n1189), .A2(n1188), .ZN(n1584) );
  NAND2_X1 U1052 ( .A1(n1230), .A2(n1229), .ZN(n1240) );
  NAND2_X1 U1053 ( .A1(n1232), .A2(n1231), .ZN(n1229) );
  NAND2_X1 U1054 ( .A1(n1234), .A2(n1228), .ZN(n1230) );
  NAND2_X1 U1055 ( .A1(n1227), .A2(n1226), .ZN(n1228) );
  OR2_X1 U1056 ( .A1(n1520), .A2(n1519), .ZN(n1525) );
  CLKBUF_X1 U1057 ( .A(n1860), .Z(n982) );
  CLKBUF_X1 U1058 ( .A(n940), .Z(n1676) );
  CLKBUF_X1 U1059 ( .A(w_to_multf[7]), .Z(n950) );
  NAND2_X1 U1060 ( .A1(n1427), .A2(n1426), .ZN(n1428) );
  NAND2_X1 U1061 ( .A1(n1195), .A2(n1196), .ZN(n957) );
  NAND2_X1 U1062 ( .A1(n1195), .A2(n1196), .ZN(n1373) );
  INV_X1 U1063 ( .A(n1232), .ZN(n1227) );
  INV_X1 U1064 ( .A(n1231), .ZN(n1226) );
  XNOR2_X1 U1065 ( .A(n1389), .B(n1388), .ZN(n1479) );
  XNOR2_X1 U1066 ( .A(n1234), .B(n1233), .ZN(n1239) );
  XNOR2_X1 U1067 ( .A(n1232), .B(n1231), .ZN(n1233) );
  INV_X1 U1068 ( .A(n978), .ZN(n1621) );
  CLKBUF_X1 U1069 ( .A(n1629), .Z(n993) );
  OAI21_X1 U1070 ( .B1(n1248), .B2(n1247), .A(n1246), .ZN(n1250) );
  XNOR2_X1 U1071 ( .A(n1175), .B(n1174), .ZN(n1180) );
  XNOR2_X1 U1072 ( .A(n1173), .B(n1172), .ZN(n1174) );
  INV_X1 U1073 ( .A(n1506), .ZN(n1515) );
  NAND2_X1 U1074 ( .A1(n1147), .A2(n1146), .ZN(n1183) );
  NAND2_X1 U1075 ( .A1(n1173), .A2(n1172), .ZN(n1146) );
  NAND2_X1 U1076 ( .A1(n1175), .A2(n1145), .ZN(n1147) );
  OR2_X1 U1077 ( .A1(n1173), .A2(n1172), .ZN(n1145) );
  NOR2_X1 U1078 ( .A1(n1839), .A2(n1837), .ZN(n1788) );
  XNOR2_X1 U1079 ( .A(n1605), .B(n1604), .ZN(n1606) );
  INV_X1 U1080 ( .A(n962), .ZN(n963) );
  CLKBUF_X1 U1081 ( .A(n1790), .Z(n981) );
  CLKBUF_X1 U1082 ( .A(n1839), .Z(n980) );
  CLKBUF_X1 U1083 ( .A(n1861), .Z(n1896) );
  CLKBUF_X1 U1084 ( .A(n1836), .Z(n997) );
  CLKBUF_X1 U1085 ( .A(n1811), .Z(n1812) );
  NAND2_X1 U1086 ( .A1(n1044), .A2(n1047), .ZN(n2094) );
  OR2_X1 U1087 ( .A1(n2055), .A2(w_write_addr_x[3]), .ZN(n2068) );
  INV_X1 U1088 ( .A(n2009), .ZN(n2010) );
  BUF_X1 U1089 ( .A(n1884), .Z(n977) );
  CLKBUF_X1 U1090 ( .A(n1900), .Z(n1000) );
  INV_X1 U1091 ( .A(n2064), .ZN(n2065) );
  INV_X1 U1092 ( .A(n2066), .ZN(n2067) );
  INV_X1 U1093 ( .A(n2085), .ZN(n2086) );
  INV_X1 U1094 ( .A(n2088), .ZN(n2089) );
  INV_X1 U1095 ( .A(n2060), .ZN(n2061) );
  INV_X1 U1096 ( .A(n2062), .ZN(n2063) );
  INV_X1 U1097 ( .A(n2080), .ZN(n2081) );
  INV_X1 U1098 ( .A(n2083), .ZN(n2084) );
  INV_X1 U1099 ( .A(n2056), .ZN(n2057) );
  INV_X1 U1100 ( .A(n2058), .ZN(n2059) );
  INV_X1 U1101 ( .A(n2074), .ZN(n2075) );
  INV_X1 U1102 ( .A(n2078), .ZN(n2079) );
  INV_X1 U1103 ( .A(n2072), .ZN(n2073) );
  INV_X1 U1104 ( .A(n2091), .ZN(n2092) );
  INV_X1 U1105 ( .A(n2095), .ZN(n2096) );
  INV_X1 U1106 ( .A(n2069), .ZN(n2070) );
  NAND2_X1 U1107 ( .A1(s_valid_x), .A2(s_ready_x), .ZN(n2009) );
  NAND2_X1 U1108 ( .A1(n1010), .A2(n1804), .ZN(n1683) );
  BUF_X1 U1109 ( .A(n1801), .Z(n940) );
  BUF_X1 U1110 ( .A(n1866), .Z(n941) );
  NAND2_X1 U1111 ( .A1(n1318), .A2(n1316), .ZN(n942) );
  NAND2_X1 U1112 ( .A1(n1318), .A2(n1316), .ZN(n1289) );
  XOR2_X1 U1113 ( .A(n994), .B(n949), .Z(n1351) );
  XOR2_X1 U1114 ( .A(n1017), .B(w_to_multf[15]), .Z(n1204) );
  BUF_X1 U1115 ( .A(n1144), .Z(n944) );
  XNOR2_X1 U1116 ( .A(n1015), .B(n968), .ZN(n1374) );
  XNOR2_X1 U1117 ( .A(n1018), .B(n2106), .ZN(n1318) );
  INV_X1 U1118 ( .A(n946), .ZN(n947) );
  INV_X1 U1119 ( .A(n994), .ZN(n948) );
  INV_X1 U1120 ( .A(w_to_multf[7]), .ZN(n949) );
  BUF_X1 U1121 ( .A(n970), .Z(n952) );
  BUF_X1 U1122 ( .A(n970), .Z(n953) );
  BUF_X2 U1123 ( .A(n970), .Z(n954) );
  XNOR2_X1 U1124 ( .A(n2378), .B(n1021), .ZN(n970) );
  INV_X1 U1125 ( .A(n964), .ZN(n956) );
  INV_X1 U1126 ( .A(n968), .ZN(n958) );
  INV_X1 U1127 ( .A(n959), .ZN(n960) );
  XNOR2_X1 U1128 ( .A(n2104), .B(w_to_multx[8]), .ZN(n1196) );
  BUF_X2 U1129 ( .A(\DP_OP_65J1_123_5677/n1044 ), .Z(n961) );
  XNOR2_X1 U1130 ( .A(w_to_multx[10]), .B(w_to_multx[9]), .ZN(n965) );
  XOR2_X1 U1131 ( .A(w_to_multf[15]), .B(n1018), .Z(n1274) );
  INV_X1 U1132 ( .A(w_to_multx[13]), .ZN(n966) );
  INV_X1 U1133 ( .A(n939), .ZN(n967) );
  XNOR2_X1 U1134 ( .A(n961), .B(w_to_multf[5]), .ZN(n1252) );
  NAND2_X1 U1135 ( .A1(n1101), .A2(n965), .ZN(n1406) );
  XNOR2_X1 U1136 ( .A(n1015), .B(w_to_multx[12]), .ZN(n1093) );
  XNOR2_X1 U1137 ( .A(n1013), .B(w_to_multx[14]), .ZN(n1096) );
  XNOR2_X2 U1138 ( .A(w_to_multx[5]), .B(w_to_multx[6]), .ZN(n974) );
  XNOR2_X1 U1139 ( .A(n1857), .B(n975), .ZN(n1890) );
  AND2_X1 U1140 ( .A1(n1856), .A2(n1855), .ZN(n975) );
  XNOR2_X1 U1141 ( .A(n1018), .B(w_to_multx[4]), .ZN(n1273) );
  OR2_X1 U1142 ( .A1(n1608), .A2(n1607), .ZN(n976) );
  OR2_X1 U1143 ( .A1(n1608), .A2(n1607), .ZN(n1595) );
  NAND2_X1 U1144 ( .A1(n1203), .A2(n1113), .ZN(n1194) );
  NOR2_X1 U1145 ( .A1(n1655), .A2(\conv/prev_output [13]), .ZN(n1869) );
  AOI21_X1 U1146 ( .B1(n1566), .B2(n1565), .A(n1564), .ZN(n1582) );
  XNOR2_X1 U1147 ( .A(n1872), .B(n983), .ZN(n1972) );
  AND2_X1 U1148 ( .A1(n1871), .A2(n1870), .ZN(n983) );
  AOI21_X1 U1149 ( .B1(n1653), .B2(n1652), .A(n1651), .ZN(n984) );
  AOI21_X1 U1150 ( .B1(n1653), .B2(n1652), .A(n1651), .ZN(n1874) );
  INV_X1 U1151 ( .A(n1878), .ZN(n985) );
  NAND2_X1 U1152 ( .A1(n1583), .A2(n1647), .ZN(n986) );
  AND2_X1 U1153 ( .A1(n989), .A2(n1525), .ZN(n987) );
  AND2_X1 U1154 ( .A1(n1526), .A2(n1525), .ZN(n1614) );
  XNOR2_X1 U1155 ( .A(n1469), .B(n1473), .ZN(n1445) );
  NAND2_X1 U1156 ( .A1(n1509), .A2(n1508), .ZN(n989) );
  INV_X1 U1157 ( .A(n1122), .ZN(n1123) );
  AND2_X1 U1158 ( .A1(n1122), .A2(n1124), .ZN(n1223) );
  OAI21_X1 U1159 ( .B1(n942), .B2(n1317), .A(n1278), .ZN(n1292) );
  OAI21_X1 U1160 ( .B1(n1289), .B2(n1118), .A(n1117), .ZN(n1122) );
  XOR2_X1 U1161 ( .A(n996), .B(n1347), .Z(n1438) );
  NAND2_X1 U1162 ( .A1(n1131), .A2(n1273), .ZN(n991) );
  NAND2_X1 U1163 ( .A1(n1131), .A2(n1273), .ZN(n1261) );
  XNOR2_X1 U1164 ( .A(n1265), .B(n1264), .ZN(n1216) );
  XNOR2_X1 U1165 ( .A(n1216), .B(n1263), .ZN(n1241) );
  XNOR2_X1 U1166 ( .A(n1609), .B(n1596), .ZN(n1597) );
  OR2_X2 U1167 ( .A1(n1005), .A2(n1006), .ZN(n2007) );
  XNOR2_X1 U1168 ( .A(n1016), .B(n995), .ZN(n1094) );
  NAND2_X1 U1169 ( .A1(n1327), .A2(n1326), .ZN(n996) );
  NAND2_X1 U1170 ( .A1(n1327), .A2(n1326), .ZN(n1628) );
  NAND2_X2 U1171 ( .A1(n1908), .A2(n1804), .ZN(n1916) );
  NAND2_X1 U1172 ( .A1(n1369), .A2(n1368), .ZN(n1370) );
  XNOR2_X1 U1173 ( .A(n1905), .B(n998), .ZN(n1978) );
  AND2_X1 U1174 ( .A1(n1904), .A2(n1903), .ZN(n998) );
  XNOR2_X1 U1175 ( .A(n1879), .B(n999), .ZN(n1975) );
  AND2_X1 U1176 ( .A1(n1878), .A2(n1877), .ZN(n999) );
  NOR2_X1 U1177 ( .A1(n1004), .A2(n1683), .ZN(\conv/N125 ) );
  XNOR2_X1 U1178 ( .A(n1863), .B(n1001), .ZN(n1981) );
  AND2_X1 U1179 ( .A1(n1862), .A2(n1895), .ZN(n1001) );
  AND3_X2 U1180 ( .A1(n1909), .A2(n1908), .A3(n1804), .ZN(n1002) );
  AND3_X2 U1181 ( .A1(n1909), .A2(n1908), .A3(n1804), .ZN(n1008) );
  NOR2_X1 U1182 ( .A1(n1482), .A2(n1481), .ZN(n1003) );
  AND2_X1 U1183 ( .A1(n1909), .A2(n1908), .ZN(n1004) );
  NAND2_X1 U1184 ( .A1(n1804), .A2(n2099), .ZN(n1006) );
  OR2_X4 U1185 ( .A1(n1005), .A2(n1006), .ZN(n1007) );
  BUF_X2 U1186 ( .A(n1845), .Z(n1900) );
  NOR2_X1 U1187 ( .A1(n1511), .A2(n1510), .ZN(n1009) );
  AND2_X1 U1188 ( .A1(n1682), .A2(n1803), .ZN(n1010) );
  XOR2_X1 U1189 ( .A(n1511), .B(n1510), .Z(n1011) );
  NOR2_X1 U1190 ( .A1(n1062), .A2(n1061), .ZN(n1012) );
  OR2_X1 U1191 ( .A1(n1472), .A2(n1471), .ZN(n1014) );
  XNOR2_X1 U1192 ( .A(n1588), .B(n1587), .ZN(n1019) );
  XOR2_X1 U1193 ( .A(n1616), .B(n1577), .Z(n1020) );
  XOR2_X1 U1194 ( .A(n1553), .B(n1566), .Z(n1023) );
  XOR2_X1 U1195 ( .A(n1513), .B(n1512), .Z(n1024) );
  XOR2_X1 U1196 ( .A(n1501), .B(n1500), .Z(n1025) );
  AND2_X1 U1197 ( .A1(n1647), .A2(n2098), .ZN(n1026) );
  XNOR2_X1 U1198 ( .A(n1463), .B(n1532), .ZN(n1027) );
  XNOR2_X1 U1199 ( .A(n1547), .B(n1551), .ZN(n1028) );
  NOR2_X1 U1200 ( .A1(n1501), .A2(n1500), .ZN(n1029) );
  NOR2_X1 U1201 ( .A1(w_to_multf[1]), .A2(n1013), .ZN(n1030) );
  XOR2_X1 U1202 ( .A(n1568), .B(n1567), .Z(n1031) );
  XOR2_X1 U1203 ( .A(n1534), .B(n1539), .Z(n1032) );
  NAND2_X1 U1204 ( .A1(n1524), .A2(n1532), .ZN(n1033) );
  NAND2_X1 U1205 ( .A1(n963), .A2(w_to_multx[0]), .ZN(n1034) );
  XNOR2_X1 U1206 ( .A(n1582), .B(n1581), .ZN(n1035) );
  NOR2_X1 U1207 ( .A1(n1072), .A2(n1071), .ZN(n1036) );
  NOR2_X1 U1208 ( .A1(n1082), .A2(n1081), .ZN(n1037) );
  NOR2_X1 U1209 ( .A1(n1092), .A2(n1091), .ZN(n1038) );
  XOR2_X1 U1210 ( .A(n1542), .B(n1545), .Z(n1040) );
  NOR2_X1 U1212 ( .A1(reset), .A2(\cx/overflow ), .ZN(s_ready_x) );
  AOI22_X1 U1213 ( .A1(n2010), .A2(w_write_addr_x[2]), .B1(w_read_addr_x[2]), 
        .B2(n2009), .ZN(n1043) );
  AOI22_X1 U1214 ( .A1(n2010), .A2(w_write_addr_x[1]), .B1(w_read_addr_x[1]), 
        .B2(n2009), .ZN(n1048) );
  NAND2_X1 U1215 ( .A1(n1043), .A2(n1048), .ZN(n2077) );
  NOR2_X1 U1216 ( .A1(n2009), .A2(n2109), .ZN(n2076) );
  AOI21_X1 U1217 ( .B1(w_read_addr_x[3]), .B2(n2009), .A(n2076), .ZN(n1041) );
  NOR2_X1 U1218 ( .A1(n2009), .A2(n2108), .ZN(n2032) );
  AOI21_X1 U1219 ( .B1(w_read_addr_x[0]), .B2(n2009), .A(n2032), .ZN(n1042) );
  NAND2_X1 U1220 ( .A1(n1041), .A2(n1042), .ZN(n1053) );
  NOR2_X2 U1221 ( .A1(n2077), .A2(n1053), .ZN(n1946) );
  INV_X1 U1222 ( .A(n1042), .ZN(n1045) );
  NAND2_X1 U1223 ( .A1(n1041), .A2(n1045), .ZN(n1054) );
  NOR2_X2 U1224 ( .A1(n2077), .A2(n1054), .ZN(n1945) );
  AOI22_X1 U1225 ( .A1(n1946), .A2(\mx/mem[0][2] ), .B1(n1945), .B2(
        \mx/mem[1][2] ), .ZN(n1052) );
  INV_X1 U1226 ( .A(n1048), .ZN(n1044) );
  INV_X1 U1227 ( .A(n1043), .ZN(n1047) );
  NOR2_X2 U1228 ( .A1(n2094), .A2(n1053), .ZN(n1948) );
  NOR2_X2 U1229 ( .A1(n2094), .A2(n1054), .ZN(n1947) );
  AOI22_X1 U1230 ( .A1(n1948), .A2(\mx/mem[6][2] ), .B1(n1947), .B2(
        \mx/mem[7][2] ), .ZN(n1051) );
  INV_X1 U1231 ( .A(n1041), .ZN(n1046) );
  NAND2_X1 U1232 ( .A1(n1042), .A2(n1046), .ZN(n1055) );
  NAND2_X1 U1233 ( .A1(n1044), .A2(n1043), .ZN(n2082) );
  NOR2_X2 U1234 ( .A1(n1055), .A2(n2082), .ZN(n1950) );
  NAND2_X1 U1235 ( .A1(n1046), .A2(n1045), .ZN(n1056) );
  NOR2_X2 U1236 ( .A1(n2082), .A2(n1056), .ZN(n1949) );
  AOI22_X1 U1237 ( .A1(n1950), .A2(\mx/mem[10][2] ), .B1(n1949), .B2(
        \mx/mem[11][2] ), .ZN(n1050) );
  NAND2_X1 U1238 ( .A1(n1048), .A2(n1047), .ZN(n2087) );
  NOR2_X2 U1239 ( .A1(n2087), .A2(n1053), .ZN(n1952) );
  NOR2_X2 U1240 ( .A1(n2087), .A2(n1054), .ZN(n1951) );
  AOI22_X1 U1241 ( .A1(n1952), .A2(\mx/mem[4][2] ), .B1(n1951), .B2(
        \mx/mem[5][2] ), .ZN(n1049) );
  NAND4_X1 U1242 ( .A1(n1052), .A2(n1051), .A3(n1050), .A4(n1049), .ZN(n1062)
         );
  NOR2_X2 U1243 ( .A1(n1055), .A2(n2077), .ZN(n1958) );
  NOR2_X2 U1244 ( .A1(n1056), .A2(n2077), .ZN(n1957) );
  AOI22_X1 U1245 ( .A1(n1958), .A2(\mx/mem[8][2] ), .B1(n1957), .B2(
        \mx/mem[9][2] ), .ZN(n1060) );
  NOR2_X2 U1246 ( .A1(n1055), .A2(n2094), .ZN(n1960) );
  NOR2_X2 U1247 ( .A1(n1056), .A2(n2094), .ZN(n1959) );
  AOI22_X1 U1248 ( .A1(n1960), .A2(\mx/mem[14][2] ), .B1(n1959), .B2(
        \mx/mem[15][2] ), .ZN(n1059) );
  NOR2_X2 U1249 ( .A1(n2082), .A2(n1053), .ZN(n1962) );
  NOR2_X2 U1250 ( .A1(n2082), .A2(n1054), .ZN(n1961) );
  AOI22_X1 U1251 ( .A1(n1962), .A2(\mx/mem[2][2] ), .B1(n1961), .B2(
        \mx/mem[3][2] ), .ZN(n1058) );
  NOR2_X2 U1252 ( .A1(n1055), .A2(n2087), .ZN(n1964) );
  NOR2_X2 U1253 ( .A1(n1056), .A2(n2087), .ZN(n1963) );
  AOI22_X1 U1254 ( .A1(n1964), .A2(\mx/mem[12][2] ), .B1(n1963), .B2(
        \mx/mem[13][2] ), .ZN(n1057) );
  NAND4_X1 U1255 ( .A1(n1060), .A2(n1059), .A3(n1058), .A4(n1057), .ZN(n1061)
         );
  AOI22_X1 U1256 ( .A1(n1946), .A2(\mx/mem[0][6] ), .B1(n1945), .B2(
        \mx/mem[1][6] ), .ZN(n1066) );
  AOI22_X1 U1257 ( .A1(n1948), .A2(\mx/mem[6][6] ), .B1(n1947), .B2(
        \mx/mem[7][6] ), .ZN(n1065) );
  AOI22_X1 U1258 ( .A1(n1950), .A2(\mx/mem[10][6] ), .B1(n1949), .B2(
        \mx/mem[11][6] ), .ZN(n1064) );
  AOI22_X1 U1259 ( .A1(n1952), .A2(\mx/mem[4][6] ), .B1(n1951), .B2(
        \mx/mem[5][6] ), .ZN(n1063) );
  NAND4_X1 U1260 ( .A1(n1066), .A2(n1065), .A3(n1064), .A4(n1063), .ZN(n1072)
         );
  AOI22_X1 U1261 ( .A1(n1958), .A2(\mx/mem[8][6] ), .B1(n1957), .B2(
        \mx/mem[9][6] ), .ZN(n1070) );
  AOI22_X1 U1262 ( .A1(n1960), .A2(\mx/mem[14][6] ), .B1(n1959), .B2(
        \mx/mem[15][6] ), .ZN(n1069) );
  AOI22_X1 U1263 ( .A1(n1962), .A2(\mx/mem[2][6] ), .B1(n1961), .B2(
        \mx/mem[3][6] ), .ZN(n1068) );
  AOI22_X1 U1264 ( .A1(n1964), .A2(\mx/mem[12][6] ), .B1(n1963), .B2(
        \mx/mem[13][6] ), .ZN(n1067) );
  NAND4_X1 U1265 ( .A1(n1070), .A2(n1069), .A3(n1068), .A4(n1067), .ZN(n1071)
         );
  AOI22_X1 U1266 ( .A1(n1946), .A2(\mx/mem[0][7] ), .B1(n1945), .B2(
        \mx/mem[1][7] ), .ZN(n1076) );
  AOI22_X1 U1267 ( .A1(n1948), .A2(\mx/mem[6][7] ), .B1(n1947), .B2(
        \mx/mem[7][7] ), .ZN(n1075) );
  AOI22_X1 U1268 ( .A1(n1950), .A2(\mx/mem[10][7] ), .B1(n1949), .B2(
        \mx/mem[11][7] ), .ZN(n1074) );
  AOI22_X1 U1269 ( .A1(n1952), .A2(\mx/mem[4][7] ), .B1(n1951), .B2(
        \mx/mem[5][7] ), .ZN(n1073) );
  NAND4_X1 U1270 ( .A1(n1076), .A2(n1075), .A3(n1074), .A4(n1073), .ZN(n1082)
         );
  AOI22_X1 U1271 ( .A1(n1958), .A2(\mx/mem[8][7] ), .B1(n1957), .B2(
        \mx/mem[9][7] ), .ZN(n1080) );
  AOI22_X1 U1272 ( .A1(n1960), .A2(\mx/mem[14][7] ), .B1(n1959), .B2(
        \mx/mem[15][7] ), .ZN(n1079) );
  AOI22_X1 U1273 ( .A1(n1962), .A2(\mx/mem[2][7] ), .B1(n1961), .B2(
        \mx/mem[3][7] ), .ZN(n1078) );
  AOI22_X1 U1274 ( .A1(n1964), .A2(\mx/mem[12][7] ), .B1(n1963), .B2(
        \mx/mem[13][7] ), .ZN(n1077) );
  NAND4_X1 U1275 ( .A1(n1080), .A2(n1079), .A3(n1078), .A4(n1077), .ZN(n1081)
         );
  AOI22_X1 U1276 ( .A1(n1946), .A2(\mx/mem[0][9] ), .B1(n1945), .B2(
        \mx/mem[1][9] ), .ZN(n1086) );
  AOI22_X1 U1277 ( .A1(n1948), .A2(\mx/mem[6][9] ), .B1(n1947), .B2(
        \mx/mem[7][9] ), .ZN(n1085) );
  AOI22_X1 U1278 ( .A1(n1950), .A2(\mx/mem[10][9] ), .B1(n1949), .B2(
        \mx/mem[11][9] ), .ZN(n1084) );
  AOI22_X1 U1279 ( .A1(n1952), .A2(\mx/mem[4][9] ), .B1(n1951), .B2(
        \mx/mem[5][9] ), .ZN(n1083) );
  NAND4_X1 U1280 ( .A1(n1086), .A2(n1085), .A3(n1084), .A4(n1083), .ZN(n1092)
         );
  AOI22_X1 U1281 ( .A1(n1958), .A2(\mx/mem[8][9] ), .B1(n1957), .B2(
        \mx/mem[9][9] ), .ZN(n1090) );
  AOI22_X1 U1282 ( .A1(n1960), .A2(\mx/mem[14][9] ), .B1(n1959), .B2(
        \mx/mem[15][9] ), .ZN(n1089) );
  AOI22_X1 U1283 ( .A1(n1962), .A2(\mx/mem[2][9] ), .B1(n1961), .B2(
        \mx/mem[3][9] ), .ZN(n1088) );
  AOI22_X1 U1284 ( .A1(n1964), .A2(\mx/mem[12][9] ), .B1(n1963), .B2(
        \mx/mem[13][9] ), .ZN(n1087) );
  NAND4_X1 U1285 ( .A1(n1090), .A2(n1089), .A3(n1088), .A4(n1087), .ZN(n1091)
         );
  XNOR2_X1 U1286 ( .A(w_to_multx[15]), .B(w_to_multf[5]), .ZN(n1419) );
  XNOR2_X1 U1287 ( .A(w_to_multx[15]), .B(n949), .ZN(n1503) );
  OAI22_X1 U1288 ( .A1(n1504), .A2(n1419), .B1(n967), .B2(n1503), .ZN(n1107)
         );
  INV_X1 U1289 ( .A(n1107), .ZN(n1432) );
  XNOR2_X1 U1290 ( .A(w_to_multx[13]), .B(n951), .ZN(n1095) );
  XNOR2_X1 U1291 ( .A(w_to_multx[13]), .B(n949), .ZN(n1399) );
  OAI22_X1 U1292 ( .A1(n1402), .A2(n1095), .B1(n1400), .B2(n1399), .ZN(n1431)
         );
  OAI22_X1 U1293 ( .A1(n1402), .A2(n1399), .B1(n1095), .B2(n1400), .ZN(n1423)
         );
  XNOR2_X1 U1294 ( .A(w_to_multx[15]), .B(w_to_multf[4]), .ZN(n1420) );
  INV_X1 U1295 ( .A(n1420), .ZN(n1099) );
  INV_X1 U1296 ( .A(n1096), .ZN(n1097) );
  NAND2_X1 U1297 ( .A1(n1097), .A2(n1505), .ZN(n1098) );
  XNOR2_X1 U1298 ( .A(w_to_multx[10]), .B(w_to_multx[9]), .ZN(n1100) );
  NAND2_X1 U1299 ( .A1(n955), .A2(n971), .ZN(n1103) );
  XNOR2_X1 U1300 ( .A(n964), .B(w_to_multf[15]), .ZN(n1403) );
  INV_X1 U1301 ( .A(n1403), .ZN(n1102) );
  NAND2_X1 U1302 ( .A1(n1103), .A2(n1102), .ZN(n1421) );
  XNOR2_X1 U1303 ( .A(w_to_multx[15]), .B(n951), .ZN(n1109) );
  OAI22_X1 U1304 ( .A1(n1504), .A2(n1503), .B1(n1109), .B2(n967), .ZN(n1108)
         );
  AOI21_X1 U1305 ( .B1(n1400), .B2(n1402), .A(n1399), .ZN(n1104) );
  INV_X1 U1306 ( .A(n1104), .ZN(n1106) );
  HA_X1 U1307 ( .A(n1511), .B(n1510), .S(n1105) );
  INV_X1 U1308 ( .A(n1105), .ZN(n1112) );
  FA_X1 U1309 ( .A(n1108), .B(n1107), .CI(n1106), .CO(n1513), .S(n1510) );
  OAI22_X1 U1310 ( .A1(n1504), .A2(n1109), .B1(n967), .B2(n1503), .ZN(n1514)
         );
  INV_X1 U1311 ( .A(n1514), .ZN(n1512) );
  HA_X1 U1312 ( .A(n1513), .B(n1512), .S(n1110) );
  INV_X1 U1313 ( .A(n1110), .ZN(n1111) );
  NOR2_X1 U1314 ( .A1(n1112), .A2(n1111), .ZN(n1461) );
  XOR2_X1 U1315 ( .A(w_to_multx[3]), .B(w_to_multx[2]), .Z(n1203) );
  XNOR2_X1 U1316 ( .A(\DP_OP_65J1_123_5677/n1047 ), .B(w_to_multx[2]), .ZN(
        n1113) );
  XNOR2_X1 U1317 ( .A(n979), .B(n951), .ZN(n1193) );
  BUF_X2 U1318 ( .A(n1113), .Z(n1206) );
  OAI22_X1 U1319 ( .A1(n1194), .A2(n1204), .B1(n1193), .B2(n1206), .ZN(n1201)
         );
  NAND2_X1 U1320 ( .A1(\DP_OP_65J1_123_5677/n1047 ), .A2(n2105), .ZN(n1160) );
  XNOR2_X1 U1321 ( .A(w_to_multf[15]), .B(n973), .ZN(n1144) );
  AOI21_X1 U1322 ( .B1(n1160), .B2(n2105), .A(n1144), .ZN(n1208) );
  XNOR2_X1 U1323 ( .A(n2378), .B(n1021), .ZN(n1195) );
  INV_X1 U1324 ( .A(n952), .ZN(n1114) );
  AND2_X1 U1325 ( .A1(w_to_multf[1]), .A2(n1114), .ZN(n1200) );
  XNOR2_X1 U1326 ( .A(w_to_multx[3]), .B(w_to_multx[4]), .ZN(n1131) );
  XNOR2_X1 U1327 ( .A(n1213), .B(n958), .ZN(n1134) );
  OAI22_X1 U1328 ( .A1(n991), .A2(n1134), .B1(n1276), .B2(n1134), .ZN(n1127)
         );
  XNOR2_X1 U1329 ( .A(n973), .B(n951), .ZN(n1119) );
  OAI22_X1 U1330 ( .A1(n1160), .A2(n1119), .B1(n944), .B2(n2105), .ZN(n1126)
         );
  XNOR2_X1 U1331 ( .A(n979), .B(w_to_multf[5]), .ZN(n1121) );
  OAI22_X1 U1332 ( .A1(n1194), .A2(n1121), .B1(n1206), .B2(n1204), .ZN(n1125)
         );
  XNOR2_X1 U1333 ( .A(\DP_OP_65J1_123_5677/n1044 ), .B(n2106), .ZN(n1316) );
  XNOR2_X1 U1334 ( .A(n961), .B(n960), .ZN(n1116) );
  XNOR2_X1 U1335 ( .A(n961), .B(w_to_multf[4]), .ZN(n1210) );
  OAI22_X1 U1336 ( .A1(n942), .A2(n1116), .B1(n974), .B2(n1210), .ZN(n1225) );
  XNOR2_X1 U1337 ( .A(n1213), .B(w_to_multf[5]), .ZN(n1199) );
  OAI22_X1 U1338 ( .A1(n991), .A2(n1134), .B1(n1199), .B2(n1259), .ZN(n1224)
         );
  OR2_X1 U1339 ( .A1(w_to_multf[1]), .A2(n969), .ZN(n1115) );
  OAI22_X1 U1340 ( .A1(n1289), .A2(n969), .B1(n1115), .B2(n974), .ZN(n1124) );
  XNOR2_X1 U1341 ( .A(n961), .B(w_to_multf[1]), .ZN(n1118) );
  OR2_X1 U1342 ( .A1(n1116), .A2(n974), .ZN(n1117) );
  OAI22_X1 U1343 ( .A1(n1160), .A2(n944), .B1(n1119), .B2(n2105), .ZN(n1138)
         );
  INV_X1 U1344 ( .A(n974), .ZN(n1120) );
  AND2_X1 U1345 ( .A1(n963), .A2(n1120), .ZN(n1137) );
  XNOR2_X1 U1346 ( .A(n979), .B(n958), .ZN(n1150) );
  OAI22_X1 U1347 ( .A1(n1194), .A2(n1150), .B1(n1121), .B2(n1206), .ZN(n1136)
         );
  XNOR2_X1 U1348 ( .A(n1124), .B(n1123), .ZN(n1129) );
  FA_X1 U1349 ( .A(n1127), .B(n1126), .CI(n1125), .CO(n1236), .S(n1128) );
  FA_X1 U1350 ( .A(n1130), .B(n1129), .CI(n1128), .CO(n1188), .S(n1187) );
  OR2_X1 U1351 ( .A1(w_to_multf[1]), .A2(n1018), .ZN(n1132) );
  OAI22_X1 U1352 ( .A1(n991), .A2(n1018), .B1(n1132), .B2(n1259), .ZN(n1143)
         );
  XNOR2_X1 U1353 ( .A(w_to_multf[1]), .B(n1213), .ZN(n1133) );
  XNOR2_X1 U1354 ( .A(n1213), .B(w_to_multf[2]), .ZN(n1135) );
  OAI22_X1 U1355 ( .A1(n991), .A2(n1133), .B1(n1259), .B2(n1135), .ZN(n1142)
         );
  OAI22_X1 U1356 ( .A1(n991), .A2(n1135), .B1(n1259), .B2(n1134), .ZN(n1140)
         );
  FA_X1 U1357 ( .A(n1138), .B(n1137), .CI(n1136), .CO(n1130), .S(n1139) );
  NOR2_X1 U1358 ( .A1(n1187), .A2(n1186), .ZN(n1578) );
  NOR2_X1 U1359 ( .A1(n1584), .A2(n1578), .ZN(n1192) );
  FA_X1 U1360 ( .A(n1141), .B(n1140), .CI(n1139), .CO(n1186), .S(n1184) );
  HA_X1 U1361 ( .A(n1143), .B(n1142), .CO(n1141), .S(n1175) );
  OAI22_X1 U1362 ( .A1(n1194), .A2(n1150), .B1(n1206), .B2(n1150), .ZN(n1173)
         );
  XNOR2_X1 U1363 ( .A(n973), .B(w_to_multf[5]), .ZN(n1148) );
  OAI22_X1 U1364 ( .A1(n1160), .A2(n1148), .B1(n944), .B2(n2105), .ZN(n1172)
         );
  NOR2_X1 U1365 ( .A1(n1184), .A2(n1183), .ZN(n1548) );
  XNOR2_X1 U1366 ( .A(n973), .B(w_to_multf[4]), .ZN(n1156) );
  OAI22_X1 U1367 ( .A1(n1160), .A2(n1156), .B1(n1148), .B2(n2105), .ZN(n1178)
         );
  INV_X1 U1368 ( .A(n1259), .ZN(n1149) );
  AND2_X1 U1369 ( .A1(n963), .A2(n1149), .ZN(n1177) );
  XNOR2_X1 U1370 ( .A(n979), .B(w_to_multf[2]), .ZN(n1151) );
  OAI22_X1 U1371 ( .A1(n1194), .A2(n1151), .B1(n1206), .B2(n1150), .ZN(n1176)
         );
  XNOR2_X1 U1372 ( .A(w_to_multf[1]), .B(n979), .ZN(n1152) );
  OAI22_X1 U1373 ( .A1(n1194), .A2(n1152), .B1(n1206), .B2(n1151), .ZN(n1154)
         );
  OAI22_X1 U1374 ( .A1(n1160), .A2(n1156), .B1(n1156), .B2(n2105), .ZN(n1153)
         );
  NOR2_X1 U1375 ( .A1(n1170), .A2(n1169), .ZN(n1536) );
  HA_X1 U1376 ( .A(n1154), .B(n1153), .CO(n1169), .S(n1166) );
  OR2_X1 U1377 ( .A1(n963), .A2(n1017), .ZN(n1155) );
  OAI22_X1 U1378 ( .A1(n1194), .A2(n1017), .B1(n1155), .B2(n1206), .ZN(n1165)
         );
  NOR2_X1 U1379 ( .A1(n1166), .A2(n1165), .ZN(n1530) );
  XNOR2_X1 U1380 ( .A(n973), .B(w_to_multf[2]), .ZN(n1159) );
  OAI22_X1 U1381 ( .A1(n1160), .A2(n1159), .B1(n1156), .B2(n2105), .ZN(n1162)
         );
  INV_X1 U1382 ( .A(n1206), .ZN(n1157) );
  AND2_X1 U1383 ( .A1(n963), .A2(n1157), .ZN(n1161) );
  NOR2_X1 U1384 ( .A1(n1162), .A2(n1161), .ZN(n1533) );
  INV_X1 U1385 ( .A(n1533), .ZN(n1462) );
  OR2_X1 U1386 ( .A1(n963), .A2(n1039), .ZN(n1158) );
  NAND2_X1 U1387 ( .A1(n1158), .A2(n1160), .ZN(n1523) );
  OAI22_X1 U1388 ( .A1(n1160), .A2(n963), .B1(n1159), .B2(n2105), .ZN(n1522)
         );
  NAND2_X1 U1389 ( .A1(n1523), .A2(n1522), .ZN(n1532) );
  INV_X1 U1390 ( .A(n1532), .ZN(n1164) );
  NAND2_X1 U1391 ( .A1(n1162), .A2(n1161), .ZN(n1531) );
  INV_X1 U1392 ( .A(n1531), .ZN(n1163) );
  AOI21_X1 U1393 ( .B1(n1462), .B2(n1164), .A(n1163), .ZN(n1167) );
  NAND2_X1 U1394 ( .A1(n1166), .A2(n1165), .ZN(n1537) );
  OAI21_X1 U1395 ( .B1(n1530), .B2(n1167), .A(n1537), .ZN(n1168) );
  INV_X1 U1396 ( .A(n1168), .ZN(n1171) );
  NAND2_X1 U1397 ( .A1(n1170), .A2(n1169), .ZN(n1543) );
  OAI21_X1 U1398 ( .B1(n1536), .B2(n1171), .A(n1543), .ZN(n1182) );
  FA_X1 U1399 ( .A(n1178), .B(n1177), .CI(n1176), .CO(n1179), .S(n1170) );
  NAND2_X1 U1400 ( .A1(n1180), .A2(n1179), .ZN(n1550) );
  INV_X1 U1401 ( .A(n1550), .ZN(n1181) );
  AOI21_X1 U1402 ( .B1(n1182), .B2(n1549), .A(n1181), .ZN(n1185) );
  NAND2_X1 U1403 ( .A1(n1184), .A2(n1183), .ZN(n1563) );
  OAI21_X1 U1404 ( .B1(n1548), .B2(n1185), .A(n1563), .ZN(n1191) );
  NAND2_X1 U1405 ( .A1(n1187), .A2(n1186), .ZN(n1579) );
  OAI21_X1 U1406 ( .B1(n1584), .B2(n1579), .A(n1585), .ZN(n1190) );
  AOI21_X1 U1407 ( .B1(n1192), .B2(n1191), .A(n1190), .ZN(n1245) );
  OAI22_X1 U1408 ( .A1(n1194), .A2(n1193), .B1(n1206), .B2(n1204), .ZN(n1212)
         );
  XNOR2_X1 U1409 ( .A(w_to_multf[1]), .B(n994), .ZN(n1198) );
  XNOR2_X1 U1410 ( .A(n994), .B(w_to_multf[2]), .ZN(n1202) );
  OR2_X1 U1411 ( .A1(n1202), .A2(n953), .ZN(n1197) );
  OAI21_X1 U1412 ( .B1(n957), .B2(n1198), .A(n1197), .ZN(n1211) );
  XNOR2_X1 U1413 ( .A(n1212), .B(n1211), .ZN(n1219) );
  OAI22_X1 U1414 ( .A1(n991), .A2(n1199), .B1(n1276), .B2(n1274), .ZN(n1218)
         );
  FA_X1 U1415 ( .A(n1200), .B(n1208), .CI(n1201), .CO(n1217), .S(n1237) );
  OAI22_X1 U1416 ( .A1(n1289), .A2(n1210), .B1(n1252), .B2(n974), .ZN(n1256)
         );
  OAI22_X1 U1417 ( .A1(n1373), .A2(n1202), .B1(n953), .B2(n1271), .ZN(n1255)
         );
  INV_X1 U1418 ( .A(n1203), .ZN(n1205) );
  AOI21_X1 U1419 ( .B1(n1206), .B2(n1205), .A(n1204), .ZN(n1207) );
  INV_X1 U1420 ( .A(n1207), .ZN(n1254) );
  INV_X1 U1421 ( .A(n1208), .ZN(n1222) );
  OR2_X1 U1422 ( .A1(w_to_multf[1]), .A2(n948), .ZN(n1209) );
  OAI22_X1 U1423 ( .A1(n1373), .A2(n948), .B1(n1209), .B2(n953), .ZN(n1221) );
  OAI22_X1 U1424 ( .A1(n942), .A2(n1210), .B1(n974), .B2(n1210), .ZN(n1220) );
  OR2_X1 U1425 ( .A1(n1212), .A2(n1211), .ZN(n1247) );
  XNOR2_X1 U1426 ( .A(n1246), .B(n1247), .ZN(n1215) );
  XNOR2_X1 U1427 ( .A(n1213), .B(n951), .ZN(n1260) );
  OAI22_X1 U1428 ( .A1(n1261), .A2(n1274), .B1(n1260), .B2(n1276), .ZN(n1258)
         );
  INV_X1 U1429 ( .A(n955), .ZN(n1214) );
  AND2_X1 U1430 ( .A1(n963), .A2(n1214), .ZN(n1257) );
  XNOR2_X1 U1431 ( .A(n1215), .B(n1248), .ZN(n1263) );
  FA_X1 U1432 ( .A(n1219), .B(n1218), .CI(n1217), .CO(n1265), .S(n1234) );
  FA_X1 U1433 ( .A(n1222), .B(n1221), .CI(n1220), .CO(n1246), .S(n1232) );
  FA_X1 U1434 ( .A(n1225), .B(n1224), .CI(n1223), .CO(n1231), .S(n1235) );
  FA_X1 U1435 ( .A(n1237), .B(n1236), .CI(n1235), .CO(n1238), .S(n1189) );
  NAND2_X1 U1436 ( .A1(n1599), .A2(n1569), .ZN(n1244) );
  NAND2_X1 U1437 ( .A1(n1239), .A2(n1238), .ZN(n1573) );
  INV_X1 U1438 ( .A(n1573), .ZN(n1242) );
  AND2_X1 U1439 ( .A1(n1241), .A2(n1240), .ZN(n1598) );
  AOI21_X1 U1440 ( .B1(n1599), .B2(n1242), .A(n1598), .ZN(n1243) );
  OAI21_X1 U1441 ( .B1(n1245), .B2(n1244), .A(n1243), .ZN(n1466) );
  NAND2_X1 U1442 ( .A1(n1248), .A2(n1247), .ZN(n1249) );
  NAND2_X1 U1443 ( .A1(n1250), .A2(n1249), .ZN(n1287) );
  OAI22_X1 U1444 ( .A1(n1373), .A2(n1271), .B1(n952), .B2(n1271), .ZN(n1284)
         );
  XNOR2_X1 U1445 ( .A(w_to_multf[15]), .B(\DP_OP_65J1_123_5677/n1044 ), .ZN(
        n1317) );
  OR2_X1 U1446 ( .A1(n1317), .A2(n1318), .ZN(n1251) );
  OAI21_X1 U1447 ( .B1(n942), .B2(n1252), .A(n1251), .ZN(n1283) );
  OR2_X1 U1448 ( .A1(w_to_multf[1]), .A2(n956), .ZN(n1253) );
  OAI22_X1 U1449 ( .A1(n971), .A2(n956), .B1(n1253), .B2(n1404), .ZN(n1282) );
  FA_X1 U1450 ( .A(n1256), .B(n1255), .CI(n1254), .CO(n1270), .S(n1264) );
  HA_X1 U1451 ( .A(n1258), .B(n1257), .CO(n1269), .S(n1248) );
  OAI22_X1 U1452 ( .A1(n1261), .A2(n1260), .B1(n1259), .B2(n1274), .ZN(n1281)
         );
  XNOR2_X1 U1453 ( .A(w_to_multf[1]), .B(n945), .ZN(n1262) );
  XNOR2_X1 U1454 ( .A(n964), .B(w_to_multf[2]), .ZN(n1272) );
  OAI22_X1 U1455 ( .A1(n971), .A2(n1262), .B1(n955), .B2(n1272), .ZN(n1280) );
  XNOR2_X1 U1456 ( .A(n1281), .B(n1280), .ZN(n1268) );
  OAI21_X1 U1457 ( .B1(n1264), .B2(n1265), .A(n1263), .ZN(n1267) );
  NAND2_X1 U1458 ( .A1(n1265), .A2(n1264), .ZN(n1266) );
  NAND2_X1 U1459 ( .A1(n1267), .A2(n1266), .ZN(n1600) );
  FA_X1 U1460 ( .A(n1268), .B(n1269), .CI(n1270), .CO(n1305), .S(n1285) );
  XNOR2_X1 U1461 ( .A(n994), .B(w_to_multf[5]), .ZN(n1301) );
  OAI22_X1 U1462 ( .A1(n957), .A2(n1271), .B1(n1301), .B2(n954), .ZN(n1296) );
  XNOR2_X1 U1463 ( .A(n964), .B(w_to_multf[4]), .ZN(n1314) );
  OAI22_X1 U1464 ( .A1(n1406), .A2(n1272), .B1(n955), .B2(n1314), .ZN(n1295)
         );
  INV_X1 U1465 ( .A(n1273), .ZN(n1275) );
  AOI21_X1 U1466 ( .B1(n1276), .B2(n1275), .A(n1274), .ZN(n1277) );
  INV_X1 U1467 ( .A(n1277), .ZN(n1294) );
  XNOR2_X1 U1468 ( .A(n961), .B(n950), .ZN(n1288) );
  OR2_X1 U1469 ( .A1(n1288), .A2(n974), .ZN(n1278) );
  INV_X1 U1470 ( .A(n1400), .ZN(n1279) );
  NAND2_X1 U1471 ( .A1(n1279), .A2(w_to_multf[1]), .ZN(n1291) );
  XNOR2_X1 U1472 ( .A(n1292), .B(n1291), .ZN(n1299) );
  OR2_X1 U1473 ( .A1(n1281), .A2(n1280), .ZN(n1298) );
  FA_X1 U1474 ( .A(n1284), .B(n1282), .CI(n1283), .CO(n1297), .S(n1286) );
  FA_X1 U1475 ( .A(n1287), .B(n1286), .CI(n1285), .CO(n1607), .S(n1601) );
  NAND2_X1 U1476 ( .A1(n1603), .A2(n976), .ZN(n1329) );
  OAI22_X1 U1477 ( .A1(n942), .A2(n1288), .B1(n974), .B2(n1317), .ZN(n1307) );
  XNOR2_X1 U1478 ( .A(w_to_multf[1]), .B(w_to_multx[13]), .ZN(n1290) );
  XNOR2_X1 U1479 ( .A(w_to_multx[13]), .B(w_to_multf[2]), .ZN(n1315) );
  OAI22_X1 U1480 ( .A1(n1402), .A2(n1290), .B1(n1400), .B2(n1315), .ZN(n1306)
         );
  XNOR2_X1 U1481 ( .A(n1307), .B(n1306), .ZN(n1313) );
  INV_X1 U1482 ( .A(n1291), .ZN(n1293) );
  AND2_X1 U1483 ( .A1(n1293), .A2(n1292), .ZN(n1312) );
  FA_X1 U1484 ( .A(n1295), .B(n1296), .CI(n1294), .CO(n1311), .S(n1304) );
  OAI22_X1 U1485 ( .A1(n1406), .A2(n1314), .B1(n955), .B2(n1314), .ZN(n1310)
         );
  OR2_X1 U1486 ( .A1(w_to_multf[1]), .A2(n966), .ZN(n1300) );
  OAI22_X1 U1487 ( .A1(n1402), .A2(n966), .B1(n1300), .B2(n1400), .ZN(n1309)
         );
  XNOR2_X1 U1488 ( .A(n994), .B(n949), .ZN(n1372) );
  OAI22_X1 U1489 ( .A1(n957), .A2(n1301), .B1(n954), .B2(n1372), .ZN(n1308) );
  XNOR2_X1 U1490 ( .A(n1325), .B(n1324), .ZN(n1302) );
  XNOR2_X1 U1491 ( .A(n1323), .B(n1302), .ZN(n1333) );
  OAI22_X1 U1492 ( .A1(n1373), .A2(n1372), .B1(n1351), .B2(n954), .ZN(n1361)
         );
  AND2_X1 U1493 ( .A1(w_to_multf[1]), .A2(n939), .ZN(n1360) );
  OR2_X1 U1494 ( .A1(n1307), .A2(n1306), .ZN(n1349) );
  FA_X1 U1495 ( .A(n1310), .B(n1309), .CI(n1308), .CO(n1348), .S(n1324) );
  FA_X1 U1496 ( .A(n1313), .B(n1312), .CI(n1311), .CO(n1346), .S(n1323) );
  XNOR2_X1 U1497 ( .A(n964), .B(n947), .ZN(n1352) );
  OAI22_X1 U1498 ( .A1(n1406), .A2(n1314), .B1(n1352), .B2(n1404), .ZN(n1359)
         );
  OAI22_X1 U1499 ( .A1(n1402), .A2(n1315), .B1(n1400), .B2(n1374), .ZN(n1358)
         );
  INV_X1 U1500 ( .A(n1316), .ZN(n1319) );
  AOI21_X1 U1501 ( .B1(n1319), .B2(n974), .A(n1317), .ZN(n1320) );
  INV_X1 U1502 ( .A(n1320), .ZN(n1357) );
  XNOR2_X1 U1503 ( .A(n1346), .B(n1345), .ZN(n1321) );
  XNOR2_X1 U1504 ( .A(n1321), .B(n1344), .ZN(n1629) );
  INV_X1 U1505 ( .A(n1629), .ZN(n1328) );
  OR2_X1 U1506 ( .A1(n1325), .A2(n1324), .ZN(n1322) );
  NAND2_X1 U1507 ( .A1(n1323), .A2(n1322), .ZN(n1327) );
  NAND2_X1 U1508 ( .A1(n1325), .A2(n1324), .ZN(n1326) );
  NAND2_X1 U1509 ( .A1(n1328), .A2(n996), .ZN(n1337) );
  NAND2_X1 U1510 ( .A1(n978), .A2(n1337), .ZN(n1339) );
  NOR2_X1 U1511 ( .A1(n1329), .A2(n1339), .ZN(n1465) );
  AND2_X1 U1512 ( .A1(n1601), .A2(n1600), .ZN(n1331) );
  AND2_X1 U1513 ( .A1(n1608), .A2(n1607), .ZN(n1330) );
  OAI21_X1 U1514 ( .B1(n1331), .B2(n1330), .A(n1595), .ZN(n1340) );
  NAND2_X1 U1515 ( .A1(n1333), .A2(n1332), .ZN(n1619) );
  INV_X1 U1516 ( .A(n1619), .ZN(n1336) );
  INV_X1 U1517 ( .A(n1628), .ZN(n1334) );
  AND2_X1 U1518 ( .A1(n1334), .A2(n1629), .ZN(n1335) );
  OAI21_X1 U1519 ( .B1(n1340), .B2(n1339), .A(n1338), .ZN(n1464) );
  AOI21_X1 U1520 ( .B1(n1466), .B2(n1465), .A(n1464), .ZN(n1459) );
  INV_X1 U1521 ( .A(n1346), .ZN(n1342) );
  INV_X1 U1522 ( .A(n1345), .ZN(n1341) );
  NAND2_X1 U1523 ( .A1(n1346), .A2(n1345), .ZN(n1384) );
  NAND2_X1 U1524 ( .A1(n1385), .A2(n1384), .ZN(n1347) );
  NAND2_X1 U1525 ( .A1(n1347), .A2(n1628), .ZN(n1366) );
  FA_X1 U1526 ( .A(n1350), .B(n1349), .CI(n1348), .CO(n1387), .S(n1344) );
  INV_X1 U1527 ( .A(n1387), .ZN(n1354) );
  OAI22_X1 U1528 ( .A1(n1351), .A2(n957), .B1(n954), .B2(n1372), .ZN(n1382) );
  OAI22_X1 U1529 ( .A1(n1406), .A2(n1352), .B1(n1404), .B2(n1403), .ZN(n1381)
         );
  OAI22_X1 U1530 ( .A1(n1402), .A2(n1374), .B1(n1400), .B2(n1374), .ZN(n1380)
         );
  INV_X1 U1531 ( .A(n1386), .ZN(n1353) );
  NAND2_X1 U1532 ( .A1(n1354), .A2(n1353), .ZN(n1363) );
  XNOR2_X1 U1533 ( .A(w_to_multf[1]), .B(w_to_multx[15]), .ZN(n1355) );
  XNOR2_X1 U1534 ( .A(w_to_multx[15]), .B(w_to_multf[2]), .ZN(n1375) );
  OAI22_X1 U1535 ( .A1(n1504), .A2(n1355), .B1(n1505), .B2(n1375), .ZN(n1379)
         );
  NAND2_X1 U1536 ( .A1(n939), .A2(n1030), .ZN(n1356) );
  OAI21_X1 U1537 ( .B1(n1504), .B2(n1013), .A(n1356), .ZN(n1378) );
  XNOR2_X1 U1538 ( .A(n1379), .B(n1378), .ZN(n1367) );
  FA_X1 U1539 ( .A(n1359), .B(n1358), .CI(n1357), .CO(n1369), .S(n1345) );
  HA_X1 U1540 ( .A(n1361), .B(n1360), .CO(n1368), .S(n1350) );
  XNOR2_X1 U1541 ( .A(n1369), .B(n1368), .ZN(n1362) );
  XNOR2_X1 U1542 ( .A(n1367), .B(n1362), .ZN(n1389) );
  NAND2_X1 U1543 ( .A1(n1363), .A2(n1389), .ZN(n1365) );
  NAND2_X1 U1544 ( .A1(n1387), .A2(n1386), .ZN(n1364) );
  NAND2_X1 U1545 ( .A1(n1365), .A2(n1364), .ZN(n1476) );
  XNOR2_X1 U1546 ( .A(n1366), .B(n1476), .ZN(n1439) );
  OAI21_X1 U1547 ( .B1(n1368), .B2(n1369), .A(n1367), .ZN(n1371) );
  NAND2_X1 U1548 ( .A1(n1371), .A2(n1370), .ZN(n1412) );
  AOI21_X1 U1549 ( .B1(n1373), .B2(n953), .A(n1372), .ZN(n1392) );
  XNOR2_X1 U1550 ( .A(w_to_multx[13]), .B(w_to_multf[5]), .ZN(n1401) );
  OAI22_X1 U1551 ( .A1(n1402), .A2(n1374), .B1(n1401), .B2(n1400), .ZN(n1395)
         );
  XNOR2_X1 U1552 ( .A(n1392), .B(n1395), .ZN(n1377) );
  OAI22_X1 U1553 ( .A1(n1504), .A2(n1375), .B1(n1505), .B2(n1420), .ZN(n1396)
         );
  INV_X1 U1554 ( .A(n1396), .ZN(n1376) );
  XNOR2_X1 U1555 ( .A(n1377), .B(n1376), .ZN(n1413) );
  XNOR2_X1 U1556 ( .A(n1412), .B(n1413), .ZN(n1383) );
  OR2_X1 U1557 ( .A1(n1379), .A2(n1378), .ZN(n1409) );
  XNOR2_X1 U1558 ( .A(n945), .B(n951), .ZN(n1405) );
  OAI22_X1 U1559 ( .A1(n971), .A2(n1403), .B1(n1405), .B2(n955), .ZN(n1408) );
  FA_X1 U1560 ( .A(n1380), .B(n1381), .CI(n1382), .CO(n1407), .S(n1386) );
  XNOR2_X1 U1561 ( .A(n1383), .B(n1411), .ZN(n1475) );
  NOR2_X1 U1562 ( .A1(n1439), .A2(n1475), .ZN(n1442) );
  NAND2_X1 U1563 ( .A1(n1385), .A2(n1384), .ZN(n1467) );
  XNOR2_X1 U1564 ( .A(n1387), .B(n1386), .ZN(n1388) );
  NOR2_X1 U1565 ( .A1(n1438), .A2(n1479), .ZN(n1390) );
  NOR2_X1 U1566 ( .A1(n1442), .A2(n1390), .ZN(n1437) );
  AND2_X1 U1567 ( .A1(n1628), .A2(n1467), .ZN(n1391) );
  AND2_X1 U1568 ( .A1(n1391), .A2(n1476), .ZN(n1446) );
  OR2_X1 U1569 ( .A1(n1396), .A2(n1395), .ZN(n1394) );
  INV_X1 U1570 ( .A(n1392), .ZN(n1393) );
  NAND2_X1 U1571 ( .A1(n1394), .A2(n1393), .ZN(n1398) );
  NAND2_X1 U1572 ( .A1(n1396), .A2(n1395), .ZN(n1397) );
  NAND2_X1 U1573 ( .A1(n1398), .A2(n1397), .ZN(n1427) );
  OAI22_X1 U1574 ( .A1(n1402), .A2(n1401), .B1(n1400), .B2(n1399), .ZN(n1418)
         );
  OAI22_X1 U1575 ( .A1(n971), .A2(n1405), .B1(n955), .B2(n1403), .ZN(n1417) );
  INV_X1 U1576 ( .A(n1422), .ZN(n1416) );
  XNOR2_X1 U1577 ( .A(n1427), .B(n1426), .ZN(n1410) );
  FA_X1 U1578 ( .A(n1409), .B(n1408), .CI(n1407), .CO(n1424), .S(n1411) );
  XNOR2_X1 U1579 ( .A(n1410), .B(n1424), .ZN(n1474) );
  OAI21_X1 U1580 ( .B1(n1413), .B2(n1412), .A(n1411), .ZN(n1415) );
  NAND2_X1 U1581 ( .A1(n1413), .A2(n1412), .ZN(n1414) );
  NAND2_X1 U1582 ( .A1(n1415), .A2(n1414), .ZN(n1473) );
  NOR2_X1 U1583 ( .A1(n1446), .A2(n1445), .ZN(n1436) );
  FA_X1 U1584 ( .A(n1418), .B(n1417), .CI(n1416), .CO(n1435), .S(n1426) );
  OAI22_X1 U1585 ( .A1(n1504), .A2(n1420), .B1(n1419), .B2(n967), .ZN(n1434)
         );
  FA_X1 U1586 ( .A(n1423), .B(n1422), .CI(n1421), .CO(n1430), .S(n1433) );
  OR2_X1 U1587 ( .A1(n1426), .A2(n1427), .ZN(n1425) );
  NAND2_X1 U1588 ( .A1(n1425), .A2(n1424), .ZN(n1429) );
  NAND2_X1 U1589 ( .A1(n1429), .A2(n1428), .ZN(n1471) );
  FA_X1 U1590 ( .A(n1432), .B(n1431), .CI(n1430), .CO(n1511), .S(n1501) );
  FA_X1 U1591 ( .A(n1435), .B(n1434), .CI(n1433), .CO(n1500), .S(n1472) );
  HA_X1 U1592 ( .A(n1501), .B(n1500), .S(n1448) );
  NAND2_X1 U1593 ( .A1(n1447), .A2(n1448), .ZN(n1454) );
  NOR2_X1 U1594 ( .A1(n1436), .A2(n1454), .ZN(n1443) );
  NAND2_X1 U1595 ( .A1(n1437), .A2(n1443), .ZN(n1458) );
  NAND2_X1 U1596 ( .A1(n1438), .A2(n1479), .ZN(n1441) );
  NAND2_X1 U1597 ( .A1(n1439), .A2(n1475), .ZN(n1440) );
  OAI21_X1 U1598 ( .B1(n1442), .B2(n1441), .A(n1440), .ZN(n1444) );
  NAND2_X1 U1599 ( .A1(n1444), .A2(n1443), .ZN(n1457) );
  NAND2_X1 U1600 ( .A1(n1446), .A2(n1445), .ZN(n1453) );
  NAND3_X1 U1601 ( .A1(n990), .A2(n1447), .A3(n1448), .ZN(n1451) );
  HA_X1 U1602 ( .A(n1472), .B(n1471), .CO(n1449), .S(n1447) );
  NAND2_X1 U1603 ( .A1(n1449), .A2(n1448), .ZN(n1450) );
  AND2_X1 U1604 ( .A1(n1451), .A2(n1450), .ZN(n1452) );
  OAI21_X1 U1605 ( .B1(n1454), .B2(n1453), .A(n1452), .ZN(n1455) );
  INV_X1 U1606 ( .A(n1455), .ZN(n1456) );
  OAI211_X1 U1607 ( .C1(n1499), .C2(n1458), .A(n1457), .B(n1456), .ZN(n1460)
         );
  NAND2_X1 U1608 ( .A1(n1460), .A2(n1461), .ZN(n1521) );
  BUF_X2 U1609 ( .A(n1521), .Z(n1646) );
  NAND2_X1 U1610 ( .A1(n1462), .A2(n1531), .ZN(n1463) );
  AOI21_X1 U1611 ( .B1(n1466), .B2(n1465), .A(n1464), .ZN(n1499) );
  XNOR2_X1 U1612 ( .A(n1475), .B(n1476), .ZN(n1482) );
  OR2_X1 U1613 ( .A1(n996), .A2(n1467), .ZN(n1481) );
  NOR2_X1 U1614 ( .A1(n1482), .A2(n1481), .ZN(n1485) );
  XNOR2_X1 U1615 ( .A(n996), .B(n1467), .ZN(n1480) );
  NOR2_X1 U1616 ( .A1(n1480), .A2(n1479), .ZN(n1468) );
  NOR2_X1 U1617 ( .A1(n1485), .A2(n1468), .ZN(n1478) );
  INV_X1 U1618 ( .A(n1473), .ZN(n1470) );
  INV_X1 U1619 ( .A(n1474), .ZN(n1469) );
  NAND2_X1 U1620 ( .A1(n1470), .A2(n1469), .ZN(n1489) );
  XNOR2_X1 U1621 ( .A(n1472), .B(n1471), .ZN(n1488) );
  OAI21_X1 U1622 ( .B1(n1489), .B2(n1488), .A(n1014), .ZN(n1493) );
  XNOR2_X1 U1623 ( .A(n1474), .B(n1473), .ZN(n1486) );
  OR2_X1 U1624 ( .A1(n1476), .A2(n1475), .ZN(n1487) );
  NOR2_X1 U1625 ( .A1(n1486), .A2(n1487), .ZN(n1477) );
  NOR2_X1 U1626 ( .A1(n1493), .A2(n1477), .ZN(n1495) );
  NAND2_X1 U1627 ( .A1(n1478), .A2(n1495), .ZN(n1498) );
  NAND2_X1 U1628 ( .A1(n1480), .A2(n1479), .ZN(n1484) );
  NAND2_X1 U1629 ( .A1(n1482), .A2(n1481), .ZN(n1483) );
  OAI21_X1 U1630 ( .B1(n1003), .B2(n1484), .A(n1483), .ZN(n1496) );
  NAND2_X1 U1631 ( .A1(n1487), .A2(n1486), .ZN(n1492) );
  AND2_X1 U1632 ( .A1(n1489), .A2(n1488), .ZN(n1490) );
  NAND2_X1 U1633 ( .A1(n1490), .A2(n1014), .ZN(n1491) );
  OAI211_X1 U1634 ( .C1(n1493), .C2(n1492), .A(n1025), .B(n1491), .ZN(n1494)
         );
  AOI21_X1 U1635 ( .B1(n1496), .B2(n1495), .A(n1494), .ZN(n1497) );
  OAI21_X1 U1636 ( .B1(n1459), .B2(n1498), .A(n1497), .ZN(n1509) );
  NOR2_X1 U1637 ( .A1(n1029), .A2(n1009), .ZN(n1502) );
  OR2_X1 U1638 ( .A1(n1513), .A2(n1512), .ZN(n1517) );
  NAND2_X1 U1639 ( .A1(n1502), .A2(n1517), .ZN(n1507) );
  AOI21_X1 U1640 ( .B1(n967), .B2(n1504), .A(n1503), .ZN(n1506) );
  NOR2_X1 U1641 ( .A1(n1515), .A2(n1514), .ZN(n1519) );
  NOR2_X1 U1642 ( .A1(n1507), .A2(n1519), .ZN(n1508) );
  NAND2_X1 U1643 ( .A1(n1509), .A2(n1508), .ZN(n1526) );
  OAI21_X1 U1644 ( .B1(n1011), .B2(n1009), .A(n1024), .ZN(n1518) );
  XNOR2_X1 U1645 ( .A(n1515), .B(n1514), .ZN(n1516) );
  AOI21_X1 U1646 ( .B1(n1518), .B2(n1517), .A(n1516), .ZN(n1520) );
  OAI21_X1 U1647 ( .B1(n1646), .B2(n1027), .A(n987), .ZN(n1528) );
  NOR2_X1 U1648 ( .A1(n1528), .A2(n2101), .ZN(n1839) );
  BUF_X2 U1649 ( .A(n1521), .Z(n1640) );
  OR2_X1 U1650 ( .A1(n1523), .A2(n1522), .ZN(n1524) );
  OAI21_X1 U1651 ( .B1(n1033), .B2(n1640), .A(n1614), .ZN(n1527) );
  NOR2_X1 U1652 ( .A1(n1527), .A2(\conv/prev_output [2]), .ZN(n1837) );
  INV_X1 U1653 ( .A(n1647), .ZN(n1913) );
  NAND2_X1 U1654 ( .A1(n1913), .A2(\conv/prev_output [0]), .ZN(n1914) );
  AND2_X2 U1655 ( .A1(n1526), .A2(n1525), .ZN(n1647) );
  OAI21_X1 U1656 ( .B1(n1646), .B2(n1034), .A(n988), .ZN(n1822) );
  NAND2_X1 U1657 ( .A1(n1822), .A2(\conv/prev_output [1]), .ZN(n1823) );
  NAND2_X1 U1658 ( .A1(n1914), .A2(n1823), .ZN(n1806) );
  NOR2_X1 U1659 ( .A1(n1528), .A2(n2101), .ZN(n1529) );
  NAND2_X1 U1660 ( .A1(n1527), .A2(\conv/prev_output [2]), .ZN(n1836) );
  NAND2_X1 U1661 ( .A1(n1528), .A2(n2101), .ZN(n1840) );
  OAI21_X1 U1662 ( .B1(n1529), .B2(n1836), .A(n1840), .ZN(n1787) );
  AOI21_X1 U1663 ( .B1(n1788), .B2(n1806), .A(n1787), .ZN(n1562) );
  INV_X1 U1664 ( .A(n1530), .ZN(n1540) );
  NAND2_X1 U1665 ( .A1(n1540), .A2(n1537), .ZN(n1534) );
  OAI21_X1 U1666 ( .B1(n1533), .B2(n1532), .A(n1531), .ZN(n1539) );
  OR2_X1 U1667 ( .A1(n1640), .A2(n1032), .ZN(n1535) );
  NAND2_X1 U1668 ( .A1(n1535), .A2(n1647), .ZN(n1556) );
  NOR2_X1 U1669 ( .A1(n1556), .A2(\conv/prev_output [4]), .ZN(n1810) );
  INV_X1 U1670 ( .A(n1536), .ZN(n1546) );
  NAND2_X1 U1671 ( .A1(n1546), .A2(n1543), .ZN(n1542) );
  INV_X1 U1672 ( .A(n1537), .ZN(n1538) );
  AOI21_X1 U1673 ( .B1(n1540), .B2(n1539), .A(n1538), .ZN(n1541) );
  INV_X1 U1674 ( .A(n1541), .ZN(n1545) );
  OR2_X1 U1675 ( .A1(n1640), .A2(n1040), .ZN(n1557) );
  NOR2_X1 U1676 ( .A1(n1810), .A2(n1785), .ZN(n1555) );
  NAND2_X1 U1677 ( .A1(n1549), .A2(n1550), .ZN(n1547) );
  INV_X1 U1678 ( .A(n1543), .ZN(n1544) );
  AOI21_X1 U1679 ( .B1(n1546), .B2(n1545), .A(n1544), .ZN(n1551) );
  OAI21_X1 U1680 ( .B1(n1646), .B2(n1028), .A(n987), .ZN(n1559) );
  NOR2_X1 U1681 ( .A1(n1559), .A2(\conv/prev_output [6]), .ZN(n1786) );
  INV_X1 U1682 ( .A(n1548), .ZN(n1565) );
  NAND2_X1 U1683 ( .A1(n1565), .A2(n1563), .ZN(n1553) );
  INV_X1 U1684 ( .A(n1549), .ZN(n1552) );
  OAI21_X1 U1685 ( .B1(n1552), .B2(n1551), .A(n1550), .ZN(n1566) );
  OAI21_X1 U1686 ( .B1(n1023), .B2(n1640), .A(n1614), .ZN(n1794) );
  NOR2_X1 U1687 ( .A1(n1794), .A2(\conv/prev_output [7]), .ZN(n1554) );
  NOR2_X1 U1688 ( .A1(n1786), .A2(n1554), .ZN(n1561) );
  NAND2_X1 U1689 ( .A1(n1555), .A2(n1561), .ZN(n1661) );
  NAND2_X1 U1690 ( .A1(n1556), .A2(\conv/prev_output [4]), .ZN(n1811) );
  NAND2_X1 U1691 ( .A1(n1557), .A2(n987), .ZN(n1558) );
  NAND2_X1 U1692 ( .A1(n1558), .A2(\conv/prev_output [5]), .ZN(n1813) );
  OAI21_X1 U1693 ( .B1(n1785), .B2(n1811), .A(n1813), .ZN(n1790) );
  NAND2_X1 U1694 ( .A1(n1559), .A2(\conv/prev_output [6]), .ZN(n1831) );
  NAND2_X1 U1695 ( .A1(n1794), .A2(\conv/prev_output [7]), .ZN(n1795) );
  OAI21_X1 U1696 ( .B1(n1554), .B2(n1831), .A(n1795), .ZN(n1560) );
  AOI21_X1 U1697 ( .B1(n1561), .B2(n1790), .A(n1560), .ZN(n1660) );
  OAI21_X1 U1698 ( .B1(n1562), .B2(n1661), .A(n1660), .ZN(n1801) );
  INV_X1 U1699 ( .A(n1563), .ZN(n1564) );
  OAI21_X1 U1700 ( .B1(n1582), .B2(n1578), .A(n1579), .ZN(n1571) );
  INV_X1 U1701 ( .A(n1571), .ZN(n1588) );
  OAI21_X1 U1702 ( .B1(n1588), .B2(n943), .A(n1585), .ZN(n1568) );
  NAND2_X1 U1703 ( .A1(n1569), .A2(n1573), .ZN(n1567) );
  OAI21_X1 U1704 ( .B1(n1646), .B2(n1031), .A(n1647), .ZN(n1644) );
  NOR2_X1 U1705 ( .A1(n1644), .A2(\conv/prev_output [10]), .ZN(n1861) );
  INV_X1 U1706 ( .A(n1569), .ZN(n1572) );
  NOR2_X1 U1707 ( .A1(n1572), .A2(n943), .ZN(n1570) );
  NAND2_X1 U1708 ( .A1(n1571), .A2(n1570), .ZN(n1576) );
  NOR2_X1 U1709 ( .A1(n1572), .A2(n1585), .ZN(n1574) );
  NOR2_X1 U1710 ( .A1(n1574), .A2(n1242), .ZN(n1575) );
  NAND2_X1 U1711 ( .A1(n1576), .A2(n1575), .ZN(n1616) );
  INV_X1 U1712 ( .A(n1598), .ZN(n1594) );
  NAND2_X1 U1713 ( .A1(n1594), .A2(n1599), .ZN(n1577) );
  OR2_X1 U1714 ( .A1(n1646), .A2(n1020), .ZN(n1902) );
  AND2_X1 U1715 ( .A1(n988), .A2(n2100), .ZN(n1901) );
  AND2_X1 U1716 ( .A1(n1902), .A2(n1901), .ZN(n1643) );
  NOR2_X1 U1717 ( .A1(n1861), .A2(n1643), .ZN(n1591) );
  INV_X1 U1718 ( .A(n1578), .ZN(n1580) );
  NAND2_X1 U1719 ( .A1(n1580), .A2(n1579), .ZN(n1581) );
  OR2_X1 U1720 ( .A1(n1640), .A2(n1035), .ZN(n1583) );
  NAND2_X1 U1721 ( .A1(n1583), .A2(n1647), .ZN(n1639) );
  NOR2_X1 U1722 ( .A1(n986), .A2(\conv/prev_output [8]), .ZN(n1860) );
  INV_X1 U1723 ( .A(n943), .ZN(n1586) );
  NAND2_X1 U1724 ( .A1(n1586), .A2(n1585), .ZN(n1587) );
  OR2_X1 U1725 ( .A1(n1019), .A2(n1640), .ZN(n1589) );
  NOR2_X1 U1726 ( .A1(n1860), .A2(n1884), .ZN(n1590) );
  NAND2_X1 U1727 ( .A1(n1591), .A2(n1590), .ZN(n1866) );
  INV_X1 U1728 ( .A(n1599), .ZN(n1592) );
  INV_X1 U1729 ( .A(n1603), .ZN(n1593) );
  NOR2_X1 U1730 ( .A1(n1592), .A2(n1593), .ZN(n1618) );
  NAND2_X1 U1731 ( .A1(n1601), .A2(n1600), .ZN(n1602) );
  OAI21_X1 U1732 ( .B1(n1594), .B2(n1593), .A(n1602), .ZN(n1623) );
  AOI21_X1 U1733 ( .B1(n1616), .B2(n1618), .A(n1623), .ZN(n1609) );
  NAND2_X1 U1734 ( .A1(n1608), .A2(n1607), .ZN(n1620) );
  NAND2_X1 U1735 ( .A1(n976), .A2(n1620), .ZN(n1596) );
  OAI21_X1 U1736 ( .B1(n1646), .B2(n1597), .A(n988), .ZN(n1655) );
  AOI21_X1 U1737 ( .B1(n1616), .B2(n1599), .A(n1598), .ZN(n1605) );
  NAND2_X1 U1738 ( .A1(n1603), .A2(n1602), .ZN(n1604) );
  OAI21_X1 U1739 ( .B1(n1646), .B2(n1606), .A(n988), .ZN(n1654) );
  NOR2_X1 U1740 ( .A1(n1654), .A2(\conv/prev_output [12]), .ZN(n1865) );
  NOR2_X1 U1741 ( .A1(n1869), .A2(n1865), .ZN(n1615) );
  NOR2_X1 U1742 ( .A1(n1608), .A2(n1607), .ZN(n1617) );
  OAI21_X1 U1743 ( .B1(n1609), .B2(n1617), .A(n1620), .ZN(n1611) );
  NAND2_X1 U1744 ( .A1(n978), .A2(n1619), .ZN(n1610) );
  XNOR2_X1 U1745 ( .A(n1611), .B(n1610), .ZN(n1613) );
  INV_X1 U1746 ( .A(n1646), .ZN(n1612) );
  NAND2_X1 U1747 ( .A1(n1613), .A2(n1612), .ZN(n1656) );
  NAND2_X1 U1748 ( .A1(n1656), .A2(n1026), .ZN(n1856) );
  NAND2_X1 U1749 ( .A1(n1615), .A2(n1856), .ZN(n1671) );
  NOR2_X1 U1750 ( .A1(n1866), .A2(n1671), .ZN(n1668) );
  NAND2_X1 U1751 ( .A1(n1801), .A2(n1668), .ZN(n1638) );
  INV_X1 U1752 ( .A(n1616), .ZN(n1627) );
  NOR2_X1 U1753 ( .A1(n1617), .A2(n1621), .ZN(n1624) );
  NAND2_X1 U1754 ( .A1(n1618), .A2(n1624), .ZN(n1626) );
  OAI21_X1 U1755 ( .B1(n1621), .B2(n1620), .A(n1619), .ZN(n1622) );
  AOI21_X1 U1756 ( .B1(n1624), .B2(n1623), .A(n1622), .ZN(n1625) );
  OAI21_X1 U1757 ( .B1(n1627), .B2(n1626), .A(n1625), .ZN(n1633) );
  OR2_X1 U1758 ( .A1(n993), .A2(n996), .ZN(n1631) );
  NAND2_X1 U1759 ( .A1(n993), .A2(n996), .ZN(n1630) );
  NAND2_X1 U1760 ( .A1(n1631), .A2(n1630), .ZN(n1632) );
  XNOR2_X1 U1761 ( .A(n1633), .B(n1632), .ZN(n1634) );
  OAI21_X1 U1762 ( .B1(n1646), .B2(n1634), .A(n1647), .ZN(n1635) );
  INV_X1 U1763 ( .A(n1635), .ZN(n1677) );
  OR2_X1 U1764 ( .A1(n1635), .A2(n2099), .ZN(n1637) );
  NAND2_X1 U1765 ( .A1(n1635), .A2(n2099), .ZN(n1636) );
  NAND2_X1 U1766 ( .A1(n1637), .A2(n1636), .ZN(n1662) );
  NAND2_X1 U1767 ( .A1(n1638), .A2(n1662), .ZN(n1667) );
  OR2_X1 U1768 ( .A1(n1646), .A2(n1019), .ZN(n1641) );
  NAND2_X1 U1769 ( .A1(n1641), .A2(n988), .ZN(n1642) );
  NAND2_X1 U1770 ( .A1(n1642), .A2(\conv/prev_output [9]), .ZN(n1885) );
  NOR2_X1 U1771 ( .A1(n1861), .A2(n1650), .ZN(n1652) );
  AND2_X1 U1772 ( .A1(n1902), .A2(n1901), .ZN(n1650) );
  NAND2_X1 U1773 ( .A1(n1644), .A2(\conv/prev_output [10]), .ZN(n1895) );
  OR2_X1 U1774 ( .A1(n1020), .A2(n2100), .ZN(n1645) );
  OR2_X1 U1775 ( .A1(n1646), .A2(n1645), .ZN(n1649) );
  OR2_X1 U1776 ( .A1(n2100), .A2(n1647), .ZN(n1648) );
  AND2_X1 U1777 ( .A1(n1649), .A2(n1648), .ZN(n1903) );
  OAI21_X1 U1778 ( .B1(n1650), .B2(n1895), .A(n1903), .ZN(n1651) );
  NAND2_X1 U1779 ( .A1(n1654), .A2(\conv/prev_output [12]), .ZN(n1877) );
  NAND2_X1 U1780 ( .A1(n1655), .A2(\conv/prev_output [13]), .ZN(n1870) );
  OAI21_X1 U1781 ( .B1(n1869), .B2(n1877), .A(n1870), .ZN(n1850) );
  NAND2_X1 U1782 ( .A1(n1656), .A2(n987), .ZN(n1657) );
  NAND2_X1 U1783 ( .A1(n1657), .A2(\conv/prev_output [14]), .ZN(n1855) );
  INV_X1 U1784 ( .A(n1855), .ZN(n1658) );
  AOI21_X1 U1785 ( .B1(n1850), .B2(n1856), .A(n1658), .ZN(n1659) );
  OAI21_X1 U1786 ( .B1(n1874), .B2(n1671), .A(n1659), .ZN(n1666) );
  OAI21_X1 U1787 ( .B1(n1789), .B2(n1661), .A(n1660), .ZN(n1845) );
  INV_X1 U1788 ( .A(n1662), .ZN(n1663) );
  NAND3_X1 U1789 ( .A1(n1845), .A2(n1668), .A3(n1663), .ZN(n1665) );
  NAND2_X1 U1790 ( .A1(n1666), .A2(n1663), .ZN(n1664) );
  OAI211_X1 U1791 ( .C1(n1667), .C2(n1666), .A(n1664), .B(n1665), .ZN(n1909)
         );
  AOI21_X1 U1792 ( .B1(n1668), .B2(n1845), .A(n2099), .ZN(n1674) );
  INV_X1 U1793 ( .A(n1856), .ZN(n1675) );
  NAND2_X1 U1794 ( .A1(n1677), .A2(n1855), .ZN(n1669) );
  AOI21_X1 U1795 ( .B1(n1856), .B2(n1850), .A(n1669), .ZN(n1670) );
  OAI21_X1 U1796 ( .B1(n984), .B2(n1671), .A(n1670), .ZN(n1672) );
  INV_X1 U1797 ( .A(n1672), .ZN(n1673) );
  NAND2_X1 U1798 ( .A1(n1674), .A2(n1673), .ZN(n1908) );
  NOR2_X1 U1799 ( .A1(n1677), .A2(n1675), .ZN(n1679) );
  NOR2_X1 U1800 ( .A1(n1869), .A2(n1865), .ZN(n1848) );
  NAND2_X1 U1801 ( .A1(n1679), .A2(n1848), .ZN(n1681) );
  NOR2_X1 U1802 ( .A1(n1681), .A2(n941), .ZN(n1800) );
  NAND2_X1 U1803 ( .A1(n1676), .A2(n1800), .ZN(n1682) );
  NOR2_X1 U1804 ( .A1(n1677), .A2(n1855), .ZN(n1678) );
  AOI21_X1 U1805 ( .B1(n1679), .B2(n1850), .A(n1678), .ZN(n1680) );
  OAI21_X1 U1806 ( .B1(n984), .B2(n1681), .A(n1680), .ZN(n1799) );
  NAND2_X1 U1807 ( .A1(w_read_addr_f[0]), .A2(w_read_addr_f[1]), .ZN(n1689) );
  INV_X1 U1808 ( .A(n1689), .ZN(n1684) );
  NAND2_X1 U1809 ( .A1(n2009), .A2(n1684), .ZN(\mf/N15 ) );
  NOR4_X1 U1810 ( .A1(\cc/hold_state ), .A2(m_valid_y), .A3(\cc/en_val_y ), 
        .A4(n2110), .ZN(n1692) );
  AOI21_X1 U1811 ( .B1(m_valid_y), .B2(m_ready_y), .A(reset), .ZN(n2021) );
  OAI21_X1 U1812 ( .B1(n1692), .B2(n2111), .A(n2021), .ZN(n928) );
  NOR2_X1 U1813 ( .A1(n2117), .A2(w_read_addr_f[0]), .ZN(n1685) );
  AND2_X1 U1814 ( .A1(n2009), .A2(n1685), .ZN(\mf/N13 ) );
  INV_X1 U1815 ( .A(\mf/N13 ), .ZN(\mf/N14 ) );
  OAI21_X1 U1816 ( .B1(w_read_addr_f[0]), .B2(w_read_addr_f[1]), .A(n1689), 
        .ZN(n1686) );
  INV_X1 U1817 ( .A(n1686), .ZN(n1687) );
  AND2_X1 U1818 ( .A1(n2009), .A2(n1687), .ZN(\mf/N17 ) );
  NAND3_X1 U1819 ( .A1(\cc/number_x [3]), .A2(\cc/number_x [0]), .A3(
        \cc/number_x [2]), .ZN(n1688) );
  NOR4_X1 U1820 ( .A1(\cc/number_x [1]), .A2(\cc/hold_state ), .A3(n1689), 
        .A4(n1688), .ZN(n2022) );
  NOR2_X1 U1821 ( .A1(reset), .A2(n2022), .ZN(n2035) );
  NOR3_X1 U1822 ( .A1(\cc/hold_state ), .A2(m_valid_y), .A3(\cc/en_val_y ), 
        .ZN(n1690) );
  NAND3_X1 U1823 ( .A1(w_read_addr_f[0]), .A2(w_read_addr_f[1]), .A3(n1690), 
        .ZN(n2044) );
  NAND2_X1 U1824 ( .A1(n2035), .A2(n2044), .ZN(n2039) );
  INV_X1 U1825 ( .A(n1692), .ZN(n2013) );
  AOI21_X1 U1826 ( .B1(w_read_addr_f[0]), .B2(n1692), .A(w_read_addr_f[1]), 
        .ZN(n1691) );
  NOR2_X1 U1827 ( .A1(n2039), .A2(n1691), .ZN(n919) );
  INV_X1 U1828 ( .A(n2039), .ZN(n2012) );
  NAND2_X1 U1829 ( .A1(n2012), .A2(n1692), .ZN(n2047) );
  NAND2_X1 U1830 ( .A1(n2012), .A2(n2013), .ZN(n2046) );
  INV_X1 U1831 ( .A(n2046), .ZN(n1693) );
  NAND2_X1 U1832 ( .A1(n1693), .A2(w_read_addr_f[0]), .ZN(n1694) );
  OAI21_X1 U1833 ( .B1(w_read_addr_f[0]), .B2(n2047), .A(n1694), .ZN(n920) );
  AOI22_X1 U1834 ( .A1(n1946), .A2(\mx/mem[0][15] ), .B1(n1945), .B2(
        \mx/mem[1][15] ), .ZN(n1698) );
  AOI22_X1 U1835 ( .A1(n1948), .A2(\mx/mem[6][15] ), .B1(n1947), .B2(
        \mx/mem[7][15] ), .ZN(n1697) );
  AOI22_X1 U1836 ( .A1(n1950), .A2(\mx/mem[10][15] ), .B1(n1949), .B2(
        \mx/mem[11][15] ), .ZN(n1696) );
  AOI22_X1 U1837 ( .A1(n1952), .A2(\mx/mem[4][15] ), .B1(n1951), .B2(
        \mx/mem[5][15] ), .ZN(n1695) );
  NAND4_X1 U1838 ( .A1(n1698), .A2(n1697), .A3(n1696), .A4(n1695), .ZN(n1704)
         );
  AOI22_X1 U1839 ( .A1(n1958), .A2(\mx/mem[8][15] ), .B1(n1957), .B2(
        \mx/mem[9][15] ), .ZN(n1702) );
  AOI22_X1 U1840 ( .A1(n1960), .A2(\mx/mem[14][15] ), .B1(n1959), .B2(
        \mx/mem[15][15] ), .ZN(n1701) );
  AOI22_X1 U1841 ( .A1(n1962), .A2(\mx/mem[2][15] ), .B1(n1961), .B2(
        \mx/mem[3][15] ), .ZN(n1700) );
  AOI22_X1 U1842 ( .A1(n1964), .A2(\mx/mem[12][15] ), .B1(n1963), .B2(
        \mx/mem[13][15] ), .ZN(n1699) );
  NAND4_X1 U1843 ( .A1(n1702), .A2(n1701), .A3(n1700), .A4(n1699), .ZN(n1703)
         );
  OR2_X1 U1844 ( .A1(n1704), .A2(n1703), .ZN(\mx/N14 ) );
  AOI22_X1 U1845 ( .A1(n1946), .A2(\mx/mem[0][4] ), .B1(n1945), .B2(
        \mx/mem[1][4] ), .ZN(n1708) );
  AOI22_X1 U1846 ( .A1(n1948), .A2(\mx/mem[6][4] ), .B1(n1947), .B2(
        \mx/mem[7][4] ), .ZN(n1707) );
  AOI22_X1 U1847 ( .A1(n1950), .A2(\mx/mem[10][4] ), .B1(n1949), .B2(
        \mx/mem[11][4] ), .ZN(n1706) );
  AOI22_X1 U1848 ( .A1(n1952), .A2(\mx/mem[4][4] ), .B1(n1951), .B2(
        \mx/mem[5][4] ), .ZN(n1705) );
  NAND4_X1 U1849 ( .A1(n1708), .A2(n1707), .A3(n1706), .A4(n1705), .ZN(n1714)
         );
  AOI22_X1 U1850 ( .A1(n1958), .A2(\mx/mem[8][4] ), .B1(n1957), .B2(
        \mx/mem[9][4] ), .ZN(n1712) );
  AOI22_X1 U1851 ( .A1(n1960), .A2(\mx/mem[14][4] ), .B1(n1959), .B2(
        \mx/mem[15][4] ), .ZN(n1711) );
  AOI22_X1 U1852 ( .A1(n1962), .A2(\mx/mem[2][4] ), .B1(n1961), .B2(
        \mx/mem[3][4] ), .ZN(n1710) );
  AOI22_X1 U1853 ( .A1(n1964), .A2(\mx/mem[12][4] ), .B1(n1963), .B2(
        \mx/mem[13][4] ), .ZN(n1709) );
  NAND4_X1 U1854 ( .A1(n1712), .A2(n1711), .A3(n1710), .A4(n1709), .ZN(n1713)
         );
  OR2_X1 U1855 ( .A1(n1714), .A2(n1713), .ZN(\mx/N25 ) );
  AOI22_X1 U1856 ( .A1(n1946), .A2(\mx/mem[0][0] ), .B1(n1945), .B2(
        \mx/mem[1][0] ), .ZN(n1718) );
  AOI22_X1 U1857 ( .A1(n1948), .A2(\mx/mem[6][0] ), .B1(n1947), .B2(
        \mx/mem[7][0] ), .ZN(n1717) );
  AOI22_X1 U1858 ( .A1(n1950), .A2(\mx/mem[10][0] ), .B1(n1949), .B2(
        \mx/mem[11][0] ), .ZN(n1716) );
  AOI22_X1 U1859 ( .A1(n1952), .A2(\mx/mem[4][0] ), .B1(n1951), .B2(
        \mx/mem[5][0] ), .ZN(n1715) );
  NAND4_X1 U1860 ( .A1(n1718), .A2(n1717), .A3(n1716), .A4(n1715), .ZN(n1724)
         );
  AOI22_X1 U1861 ( .A1(n1958), .A2(\mx/mem[8][0] ), .B1(n1957), .B2(
        \mx/mem[9][0] ), .ZN(n1722) );
  AOI22_X1 U1862 ( .A1(n1960), .A2(\mx/mem[14][0] ), .B1(n1959), .B2(
        \mx/mem[15][0] ), .ZN(n1721) );
  AOI22_X1 U1863 ( .A1(n1962), .A2(\mx/mem[2][0] ), .B1(n1961), .B2(
        \mx/mem[3][0] ), .ZN(n1720) );
  AOI22_X1 U1864 ( .A1(n1964), .A2(\mx/mem[12][0] ), .B1(n1963), .B2(
        \mx/mem[13][0] ), .ZN(n1719) );
  NAND4_X1 U1865 ( .A1(n1722), .A2(n1721), .A3(n1720), .A4(n1719), .ZN(n1723)
         );
  OR2_X1 U1866 ( .A1(n1724), .A2(n1723), .ZN(\mx/N29 ) );
  AOI22_X1 U1867 ( .A1(n1946), .A2(\mx/mem[0][10] ), .B1(n1945), .B2(
        \mx/mem[1][10] ), .ZN(n1728) );
  AOI22_X1 U1868 ( .A1(n1948), .A2(\mx/mem[6][10] ), .B1(n1947), .B2(
        \mx/mem[7][10] ), .ZN(n1727) );
  AOI22_X1 U1869 ( .A1(n1950), .A2(\mx/mem[10][10] ), .B1(n1949), .B2(
        \mx/mem[11][10] ), .ZN(n1726) );
  AOI22_X1 U1870 ( .A1(n1952), .A2(\mx/mem[4][10] ), .B1(n1951), .B2(
        \mx/mem[5][10] ), .ZN(n1725) );
  NAND4_X1 U1871 ( .A1(n1728), .A2(n1727), .A3(n1726), .A4(n1725), .ZN(n1734)
         );
  AOI22_X1 U1872 ( .A1(n1958), .A2(\mx/mem[8][10] ), .B1(n1957), .B2(
        \mx/mem[9][10] ), .ZN(n1732) );
  AOI22_X1 U1873 ( .A1(n1960), .A2(\mx/mem[14][10] ), .B1(n1959), .B2(
        \mx/mem[15][10] ), .ZN(n1731) );
  AOI22_X1 U1874 ( .A1(n1962), .A2(\mx/mem[2][10] ), .B1(n1961), .B2(
        \mx/mem[3][10] ), .ZN(n1730) );
  AOI22_X1 U1875 ( .A1(n1964), .A2(\mx/mem[12][10] ), .B1(n1963), .B2(
        \mx/mem[13][10] ), .ZN(n1729) );
  NAND4_X1 U1876 ( .A1(n1732), .A2(n1731), .A3(n1730), .A4(n1729), .ZN(n1733)
         );
  OR2_X1 U1877 ( .A1(n1734), .A2(n1733), .ZN(\mx/N19 ) );
  AOI22_X1 U1878 ( .A1(n1946), .A2(\mx/mem[0][12] ), .B1(n1945), .B2(
        \mx/mem[1][12] ), .ZN(n1738) );
  AOI22_X1 U1879 ( .A1(n1948), .A2(\mx/mem[6][12] ), .B1(n1947), .B2(
        \mx/mem[7][12] ), .ZN(n1737) );
  AOI22_X1 U1880 ( .A1(n1950), .A2(\mx/mem[10][12] ), .B1(n1949), .B2(
        \mx/mem[11][12] ), .ZN(n1736) );
  AOI22_X1 U1881 ( .A1(n1952), .A2(\mx/mem[4][12] ), .B1(n1951), .B2(
        \mx/mem[5][12] ), .ZN(n1735) );
  NAND4_X1 U1882 ( .A1(n1738), .A2(n1737), .A3(n1736), .A4(n1735), .ZN(n1744)
         );
  AOI22_X1 U1883 ( .A1(n1958), .A2(\mx/mem[8][12] ), .B1(n1957), .B2(
        \mx/mem[9][12] ), .ZN(n1742) );
  AOI22_X1 U1884 ( .A1(n1960), .A2(\mx/mem[14][12] ), .B1(n1959), .B2(
        \mx/mem[15][12] ), .ZN(n1741) );
  AOI22_X1 U1885 ( .A1(n1962), .A2(\mx/mem[2][12] ), .B1(n1961), .B2(
        \mx/mem[3][12] ), .ZN(n1740) );
  AOI22_X1 U1886 ( .A1(n1964), .A2(\mx/mem[12][12] ), .B1(n1963), .B2(
        \mx/mem[13][12] ), .ZN(n1739) );
  NAND4_X1 U1887 ( .A1(n1742), .A2(n1741), .A3(n1740), .A4(n1739), .ZN(n1743)
         );
  OR2_X1 U1888 ( .A1(n1744), .A2(n1743), .ZN(\mx/N17 ) );
  AOI22_X1 U1889 ( .A1(n1946), .A2(\mx/mem[0][14] ), .B1(n1945), .B2(
        \mx/mem[1][14] ), .ZN(n1748) );
  AOI22_X1 U1890 ( .A1(n1948), .A2(\mx/mem[6][14] ), .B1(n1947), .B2(
        \mx/mem[7][14] ), .ZN(n1747) );
  AOI22_X1 U1891 ( .A1(n1950), .A2(\mx/mem[10][14] ), .B1(n1949), .B2(
        \mx/mem[11][14] ), .ZN(n1746) );
  AOI22_X1 U1892 ( .A1(n1952), .A2(\mx/mem[4][14] ), .B1(n1951), .B2(
        \mx/mem[5][14] ), .ZN(n1745) );
  NAND4_X1 U1893 ( .A1(n1748), .A2(n1747), .A3(n1746), .A4(n1745), .ZN(n1754)
         );
  AOI22_X1 U1894 ( .A1(n1958), .A2(\mx/mem[8][14] ), .B1(n1957), .B2(
        \mx/mem[9][14] ), .ZN(n1752) );
  AOI22_X1 U1895 ( .A1(n1960), .A2(\mx/mem[14][14] ), .B1(n1959), .B2(
        \mx/mem[15][14] ), .ZN(n1751) );
  AOI22_X1 U1896 ( .A1(n1962), .A2(\mx/mem[2][14] ), .B1(n1961), .B2(
        \mx/mem[3][14] ), .ZN(n1750) );
  AOI22_X1 U1897 ( .A1(n1964), .A2(\mx/mem[12][14] ), .B1(n1963), .B2(
        \mx/mem[13][14] ), .ZN(n1749) );
  NAND4_X1 U1898 ( .A1(n1752), .A2(n1751), .A3(n1750), .A4(n1749), .ZN(n1753)
         );
  OR2_X1 U1899 ( .A1(n1754), .A2(n1753), .ZN(\mx/N15 ) );
  AOI22_X1 U1900 ( .A1(n1946), .A2(\mx/mem[0][8] ), .B1(n1945), .B2(
        \mx/mem[1][8] ), .ZN(n1758) );
  AOI22_X1 U1901 ( .A1(n1948), .A2(\mx/mem[6][8] ), .B1(n1947), .B2(
        \mx/mem[7][8] ), .ZN(n1757) );
  AOI22_X1 U1902 ( .A1(n1950), .A2(\mx/mem[10][8] ), .B1(n1949), .B2(
        \mx/mem[11][8] ), .ZN(n1756) );
  AOI22_X1 U1903 ( .A1(n1952), .A2(\mx/mem[4][8] ), .B1(n1951), .B2(
        \mx/mem[5][8] ), .ZN(n1755) );
  NAND4_X1 U1904 ( .A1(n1758), .A2(n1757), .A3(n1756), .A4(n1755), .ZN(n1764)
         );
  AOI22_X1 U1905 ( .A1(n1958), .A2(\mx/mem[8][8] ), .B1(n1957), .B2(
        \mx/mem[9][8] ), .ZN(n1762) );
  AOI22_X1 U1906 ( .A1(n1960), .A2(\mx/mem[14][8] ), .B1(n1959), .B2(
        \mx/mem[15][8] ), .ZN(n1761) );
  AOI22_X1 U1907 ( .A1(n1962), .A2(\mx/mem[2][8] ), .B1(n1961), .B2(
        \mx/mem[3][8] ), .ZN(n1760) );
  AOI22_X1 U1908 ( .A1(n1964), .A2(\mx/mem[12][8] ), .B1(n1963), .B2(
        \mx/mem[13][8] ), .ZN(n1759) );
  NAND4_X1 U1909 ( .A1(n1762), .A2(n1761), .A3(n1760), .A4(n1759), .ZN(n1763)
         );
  OR2_X1 U1910 ( .A1(n1764), .A2(n1763), .ZN(\mx/N21 ) );
  AOI22_X1 U1911 ( .A1(n1946), .A2(\mx/mem[0][13] ), .B1(n1945), .B2(
        \mx/mem[1][13] ), .ZN(n1768) );
  AOI22_X1 U1912 ( .A1(n1948), .A2(\mx/mem[6][13] ), .B1(n1947), .B2(
        \mx/mem[7][13] ), .ZN(n1767) );
  AOI22_X1 U1913 ( .A1(n1950), .A2(\mx/mem[10][13] ), .B1(n1949), .B2(
        \mx/mem[11][13] ), .ZN(n1766) );
  AOI22_X1 U1914 ( .A1(n1952), .A2(\mx/mem[4][13] ), .B1(n1951), .B2(
        \mx/mem[5][13] ), .ZN(n1765) );
  NAND4_X1 U1915 ( .A1(n1768), .A2(n1767), .A3(n1766), .A4(n1765), .ZN(n1774)
         );
  AOI22_X1 U1916 ( .A1(n1958), .A2(\mx/mem[8][13] ), .B1(n1957), .B2(
        \mx/mem[9][13] ), .ZN(n1772) );
  AOI22_X1 U1917 ( .A1(n1960), .A2(\mx/mem[14][13] ), .B1(n1959), .B2(
        \mx/mem[15][13] ), .ZN(n1771) );
  AOI22_X1 U1918 ( .A1(n1962), .A2(\mx/mem[2][13] ), .B1(n1961), .B2(
        \mx/mem[3][13] ), .ZN(n1770) );
  AOI22_X1 U1919 ( .A1(n1964), .A2(\mx/mem[12][13] ), .B1(n1963), .B2(
        \mx/mem[13][13] ), .ZN(n1769) );
  NAND4_X1 U1920 ( .A1(n1772), .A2(n1771), .A3(n1770), .A4(n1769), .ZN(n1773)
         );
  OR2_X1 U1921 ( .A1(n1774), .A2(n1773), .ZN(\mx/N16 ) );
  AOI22_X1 U1922 ( .A1(n1946), .A2(\mx/mem[0][11] ), .B1(n1945), .B2(
        \mx/mem[1][11] ), .ZN(n1778) );
  AOI22_X1 U1923 ( .A1(n1948), .A2(\mx/mem[6][11] ), .B1(n1947), .B2(
        \mx/mem[7][11] ), .ZN(n1777) );
  AOI22_X1 U1924 ( .A1(n1950), .A2(\mx/mem[10][11] ), .B1(n1949), .B2(
        \mx/mem[11][11] ), .ZN(n1776) );
  AOI22_X1 U1925 ( .A1(n1952), .A2(\mx/mem[4][11] ), .B1(n1951), .B2(
        \mx/mem[5][11] ), .ZN(n1775) );
  NAND4_X1 U1926 ( .A1(n1778), .A2(n1777), .A3(n1776), .A4(n1775), .ZN(n1784)
         );
  AOI22_X1 U1927 ( .A1(n1958), .A2(\mx/mem[8][11] ), .B1(n1957), .B2(
        \mx/mem[9][11] ), .ZN(n1782) );
  AOI22_X1 U1928 ( .A1(n1960), .A2(\mx/mem[14][11] ), .B1(n1959), .B2(
        \mx/mem[15][11] ), .ZN(n1781) );
  AOI22_X1 U1929 ( .A1(n1962), .A2(\mx/mem[2][11] ), .B1(n1961), .B2(
        \mx/mem[3][11] ), .ZN(n1780) );
  AOI22_X1 U1930 ( .A1(n1964), .A2(\mx/mem[12][11] ), .B1(n1963), .B2(
        \mx/mem[13][11] ), .ZN(n1779) );
  NAND4_X1 U1931 ( .A1(n1782), .A2(n1781), .A3(n1780), .A4(n1779), .ZN(n1783)
         );
  OR2_X1 U1932 ( .A1(n1784), .A2(n1783), .ZN(\mx/N18 ) );
  OR2_X1 U1933 ( .A1(n1810), .A2(n1785), .ZN(n1827) );
  INV_X1 U1934 ( .A(n1786), .ZN(n1832) );
  INV_X1 U1935 ( .A(n1832), .ZN(n1791) );
  NOR2_X1 U1936 ( .A1(n1827), .A2(n1791), .ZN(n1793) );
  AOI21_X1 U1937 ( .B1(n1788), .B2(n1806), .A(n1787), .ZN(n1789) );
  INV_X1 U1938 ( .A(n1789), .ZN(n1830) );
  INV_X1 U1939 ( .A(n981), .ZN(n1828) );
  OAI21_X1 U1940 ( .B1(n1828), .B2(n1791), .A(n1831), .ZN(n1792) );
  AOI21_X1 U1941 ( .B1(n1793), .B2(n1830), .A(n1792), .ZN(n1798) );
  OR2_X1 U1942 ( .A1(\conv/prev_output [7]), .A2(n1794), .ZN(n1796) );
  NAND2_X1 U1943 ( .A1(n1796), .A2(n1795), .ZN(n1797) );
  XOR2_X1 U1944 ( .A(n1798), .B(n1797), .Z(n1987) );
  INV_X1 U1945 ( .A(n1987), .ZN(n1805) );
  INV_X1 U1946 ( .A(n1799), .ZN(n1803) );
  NAND2_X1 U1947 ( .A1(n940), .A2(n1800), .ZN(n1802) );
  OAI21_X1 U1948 ( .B1(n1916), .B2(n1805), .A(n2007), .ZN(\conv/N117 ) );
  INV_X1 U1949 ( .A(n1806), .ZN(n1838) );
  INV_X1 U1950 ( .A(n1837), .ZN(n1807) );
  NAND2_X1 U1951 ( .A1(n1807), .A2(n997), .ZN(n1808) );
  XOR2_X1 U1952 ( .A(n1838), .B(n1808), .Z(n2002) );
  INV_X1 U1953 ( .A(n2002), .ZN(n1809) );
  OAI21_X1 U1954 ( .B1(n1916), .B2(n1809), .A(n2007), .ZN(\conv/N112 ) );
  INV_X1 U1955 ( .A(n1810), .ZN(n1819) );
  INV_X1 U1956 ( .A(n1812), .ZN(n1818) );
  AOI21_X1 U1957 ( .B1(n1830), .B2(n1819), .A(n1818), .ZN(n1816) );
  INV_X1 U1958 ( .A(n1785), .ZN(n1814) );
  NAND2_X1 U1959 ( .A1(n1814), .A2(n1813), .ZN(n1815) );
  XOR2_X1 U1960 ( .A(n1816), .B(n1815), .Z(n1993) );
  INV_X1 U1961 ( .A(n1993), .ZN(n1817) );
  OAI21_X1 U1962 ( .B1(n1916), .B2(n1817), .A(n1007), .ZN(\conv/N115 ) );
  NAND2_X1 U1963 ( .A1(n1819), .A2(n1812), .ZN(n1820) );
  XNOR2_X1 U1964 ( .A(n1830), .B(n1820), .ZN(n1996) );
  INV_X1 U1965 ( .A(n1996), .ZN(n1821) );
  OAI21_X1 U1966 ( .B1(n1916), .B2(n1821), .A(n1007), .ZN(\conv/N114 ) );
  OR2_X1 U1967 ( .A1(n1822), .A2(\conv/prev_output [1]), .ZN(n1824) );
  NAND2_X1 U1968 ( .A1(n1824), .A2(n1823), .ZN(n1825) );
  XOR2_X1 U1969 ( .A(n1825), .B(n1914), .Z(n2006) );
  INV_X1 U1970 ( .A(n2006), .ZN(n1826) );
  OAI21_X1 U1971 ( .B1(n1916), .B2(n1826), .A(n1007), .ZN(\conv/N111 ) );
  INV_X1 U1972 ( .A(n1827), .ZN(n1829) );
  AOI21_X1 U1973 ( .B1(n1830), .B2(n1829), .A(n981), .ZN(n1834) );
  NAND2_X1 U1974 ( .A1(n1832), .A2(n1831), .ZN(n1833) );
  XOR2_X1 U1975 ( .A(n1834), .B(n1833), .Z(n1990) );
  INV_X1 U1976 ( .A(n1990), .ZN(n1835) );
  OAI21_X1 U1977 ( .B1(n1916), .B2(n1835), .A(n1007), .ZN(\conv/N116 ) );
  OAI21_X1 U1978 ( .B1(n1838), .B2(n1837), .A(n997), .ZN(n1843) );
  INV_X1 U1979 ( .A(n980), .ZN(n1841) );
  NAND2_X1 U1980 ( .A1(n1841), .A2(n1840), .ZN(n1842) );
  XNOR2_X1 U1981 ( .A(n1843), .B(n1842), .ZN(n1999) );
  INV_X1 U1982 ( .A(n1999), .ZN(n1844) );
  OAI21_X1 U1983 ( .B1(n1916), .B2(n1844), .A(n1007), .ZN(\conv/N113 ) );
  INV_X1 U1984 ( .A(n982), .ZN(n1883) );
  NAND2_X1 U1985 ( .A1(n1883), .A2(n1881), .ZN(n1846) );
  XNOR2_X1 U1986 ( .A(n1000), .B(n1846), .ZN(n1984) );
  INV_X1 U1987 ( .A(n1984), .ZN(n1847) );
  OAI21_X1 U1988 ( .B1(n1916), .B2(n1847), .A(n1007), .ZN(\conv/N118 ) );
  INV_X1 U1989 ( .A(n941), .ZN(n1876) );
  INV_X1 U1990 ( .A(n1876), .ZN(n1849) );
  INV_X1 U1991 ( .A(n1848), .ZN(n1852) );
  NOR2_X1 U1992 ( .A1(n1849), .A2(n1852), .ZN(n1854) );
  INV_X1 U1993 ( .A(n1850), .ZN(n1851) );
  OAI21_X1 U1994 ( .B1(n984), .B2(n1852), .A(n1851), .ZN(n1853) );
  AOI21_X1 U1995 ( .B1(n1900), .B2(n1854), .A(n1853), .ZN(n1857) );
  NAND3_X1 U1996 ( .A1(n1004), .A2(n1890), .A3(n1804), .ZN(n1859) );
  NOR3_X2 U1997 ( .A1(c_acc), .A2(e_acc), .A3(reset), .ZN(n2004) );
  NAND2_X1 U1998 ( .A1(n2004), .A2(m_data_out_y[14]), .ZN(n1858) );
  NAND3_X1 U1999 ( .A1(n1859), .A2(n2007), .A3(n1858), .ZN(\conv/N146 ) );
  NOR2_X1 U2000 ( .A1(n982), .A2(n977), .ZN(n1892) );
  OAI21_X1 U2001 ( .B1(n1881), .B2(n977), .A(n1885), .ZN(n1894) );
  AOI21_X1 U2002 ( .B1(n1900), .B2(n1892), .A(n1894), .ZN(n1863) );
  INV_X1 U2003 ( .A(n1896), .ZN(n1862) );
  INV_X1 U2004 ( .A(n1981), .ZN(n1864) );
  OAI21_X1 U2005 ( .B1(n1864), .B2(n1916), .A(n2007), .ZN(\conv/N120 ) );
  INV_X1 U2006 ( .A(n1865), .ZN(n1878) );
  NOR2_X1 U2007 ( .A1(n941), .A2(n985), .ZN(n1868) );
  OAI21_X1 U2008 ( .B1(n1874), .B2(n985), .A(n1877), .ZN(n1867) );
  AOI21_X1 U2009 ( .B1(n1900), .B2(n1868), .A(n1867), .ZN(n1872) );
  INV_X1 U2010 ( .A(n1869), .ZN(n1871) );
  INV_X1 U2011 ( .A(n1972), .ZN(n1873) );
  OAI21_X1 U2012 ( .B1(n1873), .B2(n1916), .A(n2007), .ZN(\conv/N123 ) );
  INV_X1 U2013 ( .A(n984), .ZN(n1875) );
  AOI21_X1 U2014 ( .B1(n1900), .B2(n1876), .A(n1875), .ZN(n1879) );
  INV_X1 U2015 ( .A(n1975), .ZN(n1880) );
  OAI21_X1 U2016 ( .B1(n1880), .B2(n1916), .A(n2007), .ZN(\conv/N122 ) );
  INV_X1 U2017 ( .A(n1881), .ZN(n1882) );
  AOI21_X1 U2018 ( .B1(n1900), .B2(n1883), .A(n1882), .ZN(n1888) );
  INV_X1 U2019 ( .A(n977), .ZN(n1886) );
  NAND2_X1 U2020 ( .A1(n1886), .A2(n1885), .ZN(n1887) );
  XOR2_X1 U2021 ( .A(n1888), .B(n1887), .Z(n1910) );
  INV_X1 U2022 ( .A(n1910), .ZN(n1889) );
  OAI21_X1 U2023 ( .B1(n1889), .B2(n1916), .A(n2007), .ZN(\conv/N119 ) );
  INV_X1 U2024 ( .A(n1890), .ZN(n1891) );
  OAI21_X1 U2025 ( .B1(n1891), .B2(n1916), .A(n2007), .ZN(\conv/N124 ) );
  INV_X1 U2026 ( .A(n1892), .ZN(n1893) );
  NOR2_X1 U2027 ( .A1(n1893), .A2(n1896), .ZN(n1899) );
  INV_X1 U2028 ( .A(n1894), .ZN(n1897) );
  OAI21_X1 U2029 ( .B1(n1897), .B2(n1896), .A(n1895), .ZN(n1898) );
  AOI21_X1 U2030 ( .B1(n1900), .B2(n1899), .A(n1898), .ZN(n1905) );
  INV_X1 U2031 ( .A(n1643), .ZN(n1904) );
  INV_X1 U2032 ( .A(n1978), .ZN(n1906) );
  OAI21_X1 U2033 ( .B1(n1906), .B2(n1916), .A(n1007), .ZN(\conv/N121 ) );
  NAND2_X1 U2034 ( .A1(n2004), .A2(m_data_out_y[9]), .ZN(n1907) );
  AND2_X1 U2035 ( .A1(n2007), .A2(n1907), .ZN(n1912) );
  NAND2_X1 U2036 ( .A1(n1002), .A2(n1910), .ZN(n1911) );
  NAND2_X1 U2037 ( .A1(n1912), .A2(n1911), .ZN(\conv/N141 ) );
  OR2_X1 U2038 ( .A1(n1913), .A2(\conv/prev_output [0]), .ZN(n1915) );
  NAND2_X1 U2039 ( .A1(n1915), .A2(n1914), .ZN(n1917) );
  OAI21_X1 U2040 ( .B1(n1916), .B2(n1917), .A(n1007), .ZN(\conv/N110 ) );
  INV_X1 U2041 ( .A(n1917), .ZN(n1919) );
  AND2_X1 U2042 ( .A1(n2004), .A2(m_data_out_y[0]), .ZN(n1918) );
  AOI21_X1 U2043 ( .B1(n1002), .B2(n1919), .A(n1918), .ZN(n1920) );
  NAND2_X1 U2044 ( .A1(n1920), .A2(n1007), .ZN(\conv/N132 ) );
  NOR2_X1 U2045 ( .A1(m_ready_y), .A2(n2114), .ZN(n2018) );
  INV_X1 U2046 ( .A(reset), .ZN(n1921) );
  MUX2_X1 U2047 ( .A(\cc/hold_state ), .B(n2018), .S(n1921), .Z(n654) );
  NAND3_X1 U2048 ( .A1(\cc/number_x [1]), .A2(\cc/number_x [0]), .A3(n2035), 
        .ZN(n1922) );
  NOR2_X1 U2049 ( .A1(n2012), .A2(n1922), .ZN(n1924) );
  NAND4_X1 U2050 ( .A1(\cc/number_x [1]), .A2(\cc/number_x [0]), .A3(
        \cc/number_x [2]), .A4(n2035), .ZN(n2041) );
  OAI21_X1 U2051 ( .B1(n2044), .B2(n2041), .A(n2035), .ZN(n2042) );
  INV_X1 U2052 ( .A(n2042), .ZN(n1923) );
  MUX2_X1 U2053 ( .A(n1924), .B(n1923), .S(\cc/number_x [2]), .Z(n916) );
  AOI22_X1 U2054 ( .A1(n1946), .A2(\mx/mem[0][3] ), .B1(n1945), .B2(
        \mx/mem[1][3] ), .ZN(n1928) );
  AOI22_X1 U2055 ( .A1(n1948), .A2(\mx/mem[6][3] ), .B1(n1947), .B2(
        \mx/mem[7][3] ), .ZN(n1927) );
  AOI22_X1 U2056 ( .A1(n1950), .A2(\mx/mem[10][3] ), .B1(n1949), .B2(
        \mx/mem[11][3] ), .ZN(n1926) );
  AOI22_X1 U2057 ( .A1(n1952), .A2(\mx/mem[4][3] ), .B1(n1951), .B2(
        \mx/mem[5][3] ), .ZN(n1925) );
  NAND4_X1 U2058 ( .A1(n1928), .A2(n1927), .A3(n1926), .A4(n1925), .ZN(n1934)
         );
  AOI22_X1 U2059 ( .A1(n1958), .A2(\mx/mem[8][3] ), .B1(n1957), .B2(
        \mx/mem[9][3] ), .ZN(n1932) );
  AOI22_X1 U2060 ( .A1(n1960), .A2(\mx/mem[14][3] ), .B1(n1959), .B2(
        \mx/mem[15][3] ), .ZN(n1931) );
  AOI22_X1 U2061 ( .A1(n1962), .A2(\mx/mem[2][3] ), .B1(n1961), .B2(
        \mx/mem[3][3] ), .ZN(n1930) );
  AOI22_X1 U2062 ( .A1(n1964), .A2(\mx/mem[12][3] ), .B1(n1963), .B2(
        \mx/mem[13][3] ), .ZN(n1929) );
  NAND4_X1 U2063 ( .A1(n1932), .A2(n1931), .A3(n1930), .A4(n1929), .ZN(n1933)
         );
  OR2_X1 U2064 ( .A1(n1934), .A2(n1933), .ZN(\mx/N26 ) );
  AOI22_X1 U2065 ( .A1(n1946), .A2(\mx/mem[0][1] ), .B1(n1945), .B2(
        \mx/mem[1][1] ), .ZN(n1938) );
  AOI22_X1 U2066 ( .A1(n1948), .A2(\mx/mem[6][1] ), .B1(n1947), .B2(
        \mx/mem[7][1] ), .ZN(n1937) );
  AOI22_X1 U2067 ( .A1(n1950), .A2(\mx/mem[10][1] ), .B1(n1949), .B2(
        \mx/mem[11][1] ), .ZN(n1936) );
  AOI22_X1 U2068 ( .A1(n1952), .A2(\mx/mem[4][1] ), .B1(n1951), .B2(
        \mx/mem[5][1] ), .ZN(n1935) );
  NAND4_X1 U2069 ( .A1(n1938), .A2(n1937), .A3(n1936), .A4(n1935), .ZN(n1944)
         );
  AOI22_X1 U2070 ( .A1(n1958), .A2(\mx/mem[8][1] ), .B1(n1957), .B2(
        \mx/mem[9][1] ), .ZN(n1942) );
  AOI22_X1 U2071 ( .A1(n1960), .A2(\mx/mem[14][1] ), .B1(n1959), .B2(
        \mx/mem[15][1] ), .ZN(n1941) );
  AOI22_X1 U2072 ( .A1(n1962), .A2(\mx/mem[2][1] ), .B1(n1961), .B2(
        \mx/mem[3][1] ), .ZN(n1940) );
  AOI22_X1 U2073 ( .A1(n1964), .A2(\mx/mem[12][1] ), .B1(n1963), .B2(
        \mx/mem[13][1] ), .ZN(n1939) );
  NAND4_X1 U2074 ( .A1(n1942), .A2(n1941), .A3(n1940), .A4(n1939), .ZN(n1943)
         );
  OR2_X1 U2075 ( .A1(n1944), .A2(n1943), .ZN(\mx/N28 ) );
  AOI22_X1 U2076 ( .A1(n1946), .A2(\mx/mem[0][5] ), .B1(n1945), .B2(
        \mx/mem[1][5] ), .ZN(n1956) );
  AOI22_X1 U2077 ( .A1(n1948), .A2(\mx/mem[6][5] ), .B1(n1947), .B2(
        \mx/mem[7][5] ), .ZN(n1955) );
  AOI22_X1 U2078 ( .A1(n1950), .A2(\mx/mem[10][5] ), .B1(n1949), .B2(
        \mx/mem[11][5] ), .ZN(n1954) );
  AOI22_X1 U2079 ( .A1(n1952), .A2(\mx/mem[4][5] ), .B1(n1951), .B2(
        \mx/mem[5][5] ), .ZN(n1953) );
  NAND4_X1 U2080 ( .A1(n1956), .A2(n1955), .A3(n1954), .A4(n1953), .ZN(n1970)
         );
  AOI22_X1 U2081 ( .A1(n1958), .A2(\mx/mem[8][5] ), .B1(n1957), .B2(
        \mx/mem[9][5] ), .ZN(n1968) );
  AOI22_X1 U2082 ( .A1(n1960), .A2(\mx/mem[14][5] ), .B1(n1959), .B2(
        \mx/mem[15][5] ), .ZN(n1967) );
  AOI22_X1 U2083 ( .A1(n1962), .A2(\mx/mem[2][5] ), .B1(n1961), .B2(
        \mx/mem[3][5] ), .ZN(n1966) );
  AOI22_X1 U2084 ( .A1(n1964), .A2(\mx/mem[12][5] ), .B1(n1963), .B2(
        \mx/mem[13][5] ), .ZN(n1965) );
  NAND4_X1 U2085 ( .A1(n1968), .A2(n1967), .A3(n1966), .A4(n1965), .ZN(n1969)
         );
  OR2_X1 U2086 ( .A1(n1970), .A2(n1969), .ZN(\mx/N24 ) );
  AND2_X1 U2087 ( .A1(n2004), .A2(m_data_out_y[13]), .ZN(n1971) );
  AOI21_X1 U2088 ( .B1(n1002), .B2(n1972), .A(n1971), .ZN(n1973) );
  NAND2_X1 U2089 ( .A1(n1973), .A2(n1007), .ZN(\conv/N145 ) );
  AND2_X1 U2090 ( .A1(n2004), .A2(m_data_out_y[12]), .ZN(n1974) );
  AOI21_X1 U2091 ( .B1(n1008), .B2(n1975), .A(n1974), .ZN(n1976) );
  NAND2_X1 U2092 ( .A1(n1976), .A2(n1007), .ZN(\conv/N144 ) );
  AND2_X1 U2093 ( .A1(n2004), .A2(m_data_out_y[11]), .ZN(n1977) );
  AOI21_X1 U2094 ( .B1(n1002), .B2(n1978), .A(n1977), .ZN(n1979) );
  NAND2_X1 U2095 ( .A1(n1979), .A2(n1007), .ZN(\conv/N143 ) );
  AND2_X1 U2096 ( .A1(n2004), .A2(m_data_out_y[10]), .ZN(n1980) );
  AOI21_X1 U2097 ( .B1(n1002), .B2(n1981), .A(n1980), .ZN(n1982) );
  NAND2_X1 U2098 ( .A1(n1982), .A2(n1007), .ZN(\conv/N142 ) );
  AND2_X1 U2099 ( .A1(n2004), .A2(m_data_out_y[8]), .ZN(n1983) );
  AOI21_X1 U2100 ( .B1(n1008), .B2(n1984), .A(n1983), .ZN(n1985) );
  NAND2_X1 U2101 ( .A1(n1985), .A2(n1007), .ZN(\conv/N140 ) );
  AND2_X1 U2102 ( .A1(n2004), .A2(m_data_out_y[7]), .ZN(n1986) );
  AOI21_X1 U2103 ( .B1(n1002), .B2(n1987), .A(n1986), .ZN(n1988) );
  NAND2_X1 U2104 ( .A1(n1988), .A2(n1007), .ZN(\conv/N139 ) );
  AND2_X1 U2105 ( .A1(n2004), .A2(m_data_out_y[6]), .ZN(n1989) );
  AOI21_X1 U2106 ( .B1(n1008), .B2(n1990), .A(n1989), .ZN(n1991) );
  NAND2_X1 U2107 ( .A1(n1991), .A2(n1007), .ZN(\conv/N138 ) );
  AND2_X1 U2108 ( .A1(n2004), .A2(m_data_out_y[5]), .ZN(n1992) );
  AOI21_X1 U2109 ( .B1(n1008), .B2(n1993), .A(n1992), .ZN(n1994) );
  NAND2_X1 U2110 ( .A1(n1994), .A2(n1007), .ZN(\conv/N137 ) );
  AND2_X1 U2111 ( .A1(n2004), .A2(m_data_out_y[4]), .ZN(n1995) );
  AOI21_X1 U2112 ( .B1(n1002), .B2(n1996), .A(n1995), .ZN(n1997) );
  NAND2_X1 U2113 ( .A1(n1997), .A2(n1007), .ZN(\conv/N136 ) );
  AND2_X1 U2114 ( .A1(n2004), .A2(m_data_out_y[3]), .ZN(n1998) );
  AOI21_X1 U2115 ( .B1(n1008), .B2(n1999), .A(n1998), .ZN(n2000) );
  NAND2_X1 U2116 ( .A1(n2000), .A2(n1007), .ZN(\conv/N135 ) );
  AND2_X1 U2117 ( .A1(n2004), .A2(m_data_out_y[2]), .ZN(n2001) );
  AOI21_X1 U2118 ( .B1(n1008), .B2(n2002), .A(n2001), .ZN(n2003) );
  NAND2_X1 U2119 ( .A1(n2003), .A2(n1007), .ZN(\conv/N134 ) );
  AND2_X1 U2120 ( .A1(n2004), .A2(m_data_out_y[1]), .ZN(n2005) );
  AOI21_X1 U2121 ( .B1(n1008), .B2(n2006), .A(n2005), .ZN(n2008) );
  NAND2_X1 U2122 ( .A1(n2008), .A2(n1007), .ZN(\conv/N133 ) );
  NAND3_X1 U2123 ( .A1(n2009), .A2(w_read_addr_f[0]), .A3(n2117), .ZN(\mf/N12 ) );
  NAND2_X1 U2125 ( .A1(n2108), .A2(n2010), .ZN(n2055) );
  AOI21_X1 U2126 ( .B1(w_conv_done), .B2(n2114), .A(reset), .ZN(n2027) );
  NAND2_X1 U2127 ( .A1(n2027), .A2(n2009), .ZN(n2031) );
  NAND2_X1 U2128 ( .A1(n2055), .A2(n2031), .ZN(n2033) );
  AOI21_X1 U2129 ( .B1(n2010), .B2(n2107), .A(n2033), .ZN(n2026) );
  NAND2_X1 U2130 ( .A1(n2032), .A2(w_write_addr_x[1]), .ZN(n2011) );
  AOI22_X1 U2131 ( .A1(w_write_addr_x[2]), .A2(n2026), .B1(n2011), .B2(n2112), 
        .ZN(n921) );
  NAND2_X1 U2132 ( .A1(\cc/number_x [3]), .A2(n2035), .ZN(n2038) );
  OAI21_X1 U2133 ( .B1(n2113), .B2(n2013), .A(n2012), .ZN(n2050) );
  OAI21_X1 U2134 ( .B1(n2039), .B2(w_read_addr_x[1]), .A(n2050), .ZN(n2014) );
  INV_X1 U2135 ( .A(n2014), .ZN(n2053) );
  OAI21_X1 U2136 ( .B1(w_read_addr_x[2]), .B2(n2039), .A(n2053), .ZN(n2016) );
  NOR2_X1 U2137 ( .A1(n2113), .A2(n2047), .ZN(n2048) );
  NAND2_X1 U2138 ( .A1(w_read_addr_x[1]), .A2(n2048), .ZN(n2054) );
  NOR2_X1 U2139 ( .A1(w_read_addr_x[3]), .A2(n2054), .ZN(n2015) );
  AOI22_X1 U2140 ( .A1(w_read_addr_x[3]), .A2(n2016), .B1(w_read_addr_x[2]), 
        .B2(n2015), .ZN(n2017) );
  OAI21_X1 U2141 ( .B1(n2044), .B2(n2038), .A(n2017), .ZN(n911) );
  NOR3_X1 U2142 ( .A1(\cc/en_val_y ), .A2(reset), .A3(n2018), .ZN(\cc/N56 ) );
  NOR2_X1 U2143 ( .A1(reset), .A2(n2044), .ZN(n929) );
  NOR2_X1 U2144 ( .A1(m_valid_y), .A2(\cc/en_val_y ), .ZN(n2020) );
  INV_X1 U2145 ( .A(n2021), .ZN(n2019) );
  NOR2_X1 U2146 ( .A1(n2020), .A2(n2019), .ZN(n927) );
  OAI21_X1 U2147 ( .B1(n2022), .B2(w_conv_done), .A(n2021), .ZN(n2023) );
  INV_X1 U2148 ( .A(n2023), .ZN(n926) );
  NAND2_X1 U2149 ( .A1(n2032), .A2(n2109), .ZN(n2071) );
  INV_X1 U2150 ( .A(n2071), .ZN(n2024) );
  NOR2_X1 U2151 ( .A1(n2107), .A2(n2112), .ZN(n2028) );
  AOI22_X1 U2152 ( .A1(n2076), .A2(n2112), .B1(n2024), .B2(n2028), .ZN(n2025)
         );
  OAI21_X1 U2153 ( .B1(n2026), .B2(n2109), .A(n2025), .ZN(n925) );
  INV_X1 U2154 ( .A(n2027), .ZN(n2030) );
  NAND3_X1 U2155 ( .A1(w_write_addr_x[3]), .A2(n2032), .A3(n2028), .ZN(n2029)
         );
  OAI21_X1 U2156 ( .B1(n2030), .B2(n2110), .A(n2029), .ZN(n924) );
  OAI21_X1 U2157 ( .B1(n2108), .B2(n2031), .A(n2055), .ZN(n923) );
  OAI22_X1 U2158 ( .A1(n2107), .A2(n2033), .B1(n2032), .B2(w_write_addr_x[1]), 
        .ZN(n2121) );
  INV_X1 U2159 ( .A(n2044), .ZN(n2034) );
  OAI221_X1 U2160 ( .B1(n2034), .B2(n2115), .C1(n2044), .C2(\cc/number_x [0]), 
        .A(n2035), .ZN(n918) );
  NOR2_X1 U2161 ( .A1(n2044), .A2(n2115), .ZN(n2037) );
  INV_X1 U2162 ( .A(n2037), .ZN(n2036) );
  INV_X1 U2163 ( .A(n2035), .ZN(n2043) );
  AOI221_X1 U2164 ( .B1(\cc/number_x [1]), .B2(n2037), .C1(n2118), .C2(n2036), 
        .A(n2043), .ZN(n917) );
  NAND2_X1 U2165 ( .A1(n2039), .A2(n2038), .ZN(n2040) );
  OAI22_X1 U2166 ( .A1(n2042), .A2(n2120), .B1(n2041), .B2(n2040), .ZN(n915)
         );
  NOR2_X1 U2167 ( .A1(n2044), .A2(n2043), .ZN(n2051) );
  NAND2_X1 U2168 ( .A1(\cc/number_x [0]), .A2(n2051), .ZN(n2045) );
  OAI221_X1 U2169 ( .B1(w_read_addr_x[0]), .B2(n2047), .C1(n2113), .C2(n2046), 
        .A(n2045), .ZN(n914) );
  AOI22_X1 U2170 ( .A1(n2051), .A2(\cc/number_x [1]), .B1(n2048), .B2(n2116), 
        .ZN(n2049) );
  OAI21_X1 U2171 ( .B1(n2050), .B2(n2116), .A(n2049), .ZN(n913) );
  NAND2_X1 U2172 ( .A1(\cc/number_x [2]), .A2(n2051), .ZN(n2052) );
  OAI221_X1 U2173 ( .B1(w_read_addr_x[2]), .B2(n2054), .C1(n2119), .C2(n2053), 
        .A(n2052), .ZN(n912) );
  NOR2_X2 U2174 ( .A1(n2077), .A2(n2068), .ZN(n2056) );
  OAI22_X1 U2175 ( .A1(n2057), .A2(s_data_in_x[0]), .B1(\mx/mem[0][0] ), .B2(
        n2056), .ZN(n2122) );
  OAI22_X1 U2176 ( .A1(n2057), .A2(s_data_in_x[1]), .B1(\mx/mem[0][1] ), .B2(
        n2056), .ZN(n2123) );
  OAI22_X1 U2177 ( .A1(n2057), .A2(s_data_in_x[2]), .B1(\mx/mem[0][2] ), .B2(
        n2056), .ZN(n2124) );
  OAI22_X1 U2178 ( .A1(n2057), .A2(s_data_in_x[3]), .B1(\mx/mem[0][3] ), .B2(
        n2056), .ZN(n2125) );
  OAI22_X1 U2179 ( .A1(n2057), .A2(s_data_in_x[4]), .B1(\mx/mem[0][4] ), .B2(
        n2056), .ZN(n2126) );
  OAI22_X1 U2180 ( .A1(n2057), .A2(s_data_in_x[5]), .B1(\mx/mem[0][5] ), .B2(
        n2056), .ZN(n2127) );
  OAI22_X1 U2181 ( .A1(n2057), .A2(s_data_in_x[6]), .B1(\mx/mem[0][6] ), .B2(
        n2056), .ZN(n2128) );
  OAI22_X1 U2182 ( .A1(n2057), .A2(s_data_in_x[7]), .B1(\mx/mem[0][7] ), .B2(
        n2056), .ZN(n2129) );
  OAI22_X1 U2183 ( .A1(n2057), .A2(s_data_in_x[8]), .B1(\mx/mem[0][8] ), .B2(
        n2056), .ZN(n2130) );
  OAI22_X1 U2184 ( .A1(n2057), .A2(s_data_in_x[9]), .B1(\mx/mem[0][9] ), .B2(
        n2056), .ZN(n2131) );
  OAI22_X1 U2185 ( .A1(n2057), .A2(s_data_in_x[10]), .B1(\mx/mem[0][10] ), 
        .B2(n2056), .ZN(n2132) );
  OAI22_X1 U2186 ( .A1(n2057), .A2(s_data_in_x[11]), .B1(\mx/mem[0][11] ), 
        .B2(n2056), .ZN(n2133) );
  OAI22_X1 U2187 ( .A1(n2057), .A2(s_data_in_x[12]), .B1(\mx/mem[0][12] ), 
        .B2(n2056), .ZN(n2134) );
  OAI22_X1 U2188 ( .A1(n2057), .A2(s_data_in_x[13]), .B1(\mx/mem[0][13] ), 
        .B2(n2056), .ZN(n2135) );
  OAI22_X1 U2189 ( .A1(n2057), .A2(s_data_in_x[14]), .B1(\mx/mem[0][14] ), 
        .B2(n2056), .ZN(n2136) );
  OAI22_X1 U2190 ( .A1(n2057), .A2(s_data_in_x[15]), .B1(\mx/mem[0][15] ), 
        .B2(n2056), .ZN(n2137) );
  NOR2_X2 U2191 ( .A1(n2077), .A2(n2071), .ZN(n2058) );
  OAI22_X1 U2192 ( .A1(n2059), .A2(s_data_in_x[0]), .B1(\mx/mem[1][0] ), .B2(
        n2058), .ZN(n2138) );
  OAI22_X1 U2193 ( .A1(n2059), .A2(s_data_in_x[1]), .B1(\mx/mem[1][1] ), .B2(
        n2058), .ZN(n2139) );
  OAI22_X1 U2194 ( .A1(n2059), .A2(s_data_in_x[2]), .B1(\mx/mem[1][2] ), .B2(
        n2058), .ZN(n2140) );
  OAI22_X1 U2195 ( .A1(n2059), .A2(s_data_in_x[3]), .B1(\mx/mem[1][3] ), .B2(
        n2058), .ZN(n2141) );
  OAI22_X1 U2196 ( .A1(n2059), .A2(s_data_in_x[4]), .B1(\mx/mem[1][4] ), .B2(
        n2058), .ZN(n2142) );
  OAI22_X1 U2197 ( .A1(n2059), .A2(s_data_in_x[5]), .B1(\mx/mem[1][5] ), .B2(
        n2058), .ZN(n2143) );
  OAI22_X1 U2198 ( .A1(n2059), .A2(s_data_in_x[6]), .B1(\mx/mem[1][6] ), .B2(
        n2058), .ZN(n2144) );
  OAI22_X1 U2199 ( .A1(n2059), .A2(s_data_in_x[7]), .B1(\mx/mem[1][7] ), .B2(
        n2058), .ZN(n2145) );
  OAI22_X1 U2200 ( .A1(n2059), .A2(s_data_in_x[8]), .B1(\mx/mem[1][8] ), .B2(
        n2058), .ZN(n2146) );
  OAI22_X1 U2201 ( .A1(n2059), .A2(s_data_in_x[9]), .B1(\mx/mem[1][9] ), .B2(
        n2058), .ZN(n2147) );
  OAI22_X1 U2202 ( .A1(n2059), .A2(s_data_in_x[10]), .B1(\mx/mem[1][10] ), 
        .B2(n2058), .ZN(n2148) );
  OAI22_X1 U2203 ( .A1(n2059), .A2(s_data_in_x[11]), .B1(\mx/mem[1][11] ), 
        .B2(n2058), .ZN(n2149) );
  OAI22_X1 U2204 ( .A1(n2059), .A2(s_data_in_x[12]), .B1(\mx/mem[1][12] ), 
        .B2(n2058), .ZN(n2150) );
  OAI22_X1 U2205 ( .A1(n2059), .A2(s_data_in_x[13]), .B1(\mx/mem[1][13] ), 
        .B2(n2058), .ZN(n2151) );
  OAI22_X1 U2206 ( .A1(n2059), .A2(s_data_in_x[14]), .B1(\mx/mem[1][14] ), 
        .B2(n2058), .ZN(n2152) );
  OAI22_X1 U2207 ( .A1(n2059), .A2(s_data_in_x[15]), .B1(\mx/mem[1][15] ), 
        .B2(n2058), .ZN(n2153) );
  NOR2_X2 U2208 ( .A1(n2082), .A2(n2068), .ZN(n2060) );
  OAI22_X1 U2209 ( .A1(n2061), .A2(s_data_in_x[0]), .B1(\mx/mem[2][0] ), .B2(
        n2060), .ZN(n2154) );
  OAI22_X1 U2210 ( .A1(n2061), .A2(s_data_in_x[1]), .B1(\mx/mem[2][1] ), .B2(
        n2060), .ZN(n2155) );
  OAI22_X1 U2211 ( .A1(n2061), .A2(s_data_in_x[2]), .B1(\mx/mem[2][2] ), .B2(
        n2060), .ZN(n2156) );
  OAI22_X1 U2212 ( .A1(n2061), .A2(s_data_in_x[3]), .B1(\mx/mem[2][3] ), .B2(
        n2060), .ZN(n2157) );
  OAI22_X1 U2213 ( .A1(n2061), .A2(s_data_in_x[4]), .B1(\mx/mem[2][4] ), .B2(
        n2060), .ZN(n2158) );
  OAI22_X1 U2214 ( .A1(n2061), .A2(s_data_in_x[5]), .B1(\mx/mem[2][5] ), .B2(
        n2060), .ZN(n2159) );
  OAI22_X1 U2215 ( .A1(n2061), .A2(s_data_in_x[6]), .B1(\mx/mem[2][6] ), .B2(
        n2060), .ZN(n2160) );
  OAI22_X1 U2216 ( .A1(n2061), .A2(s_data_in_x[7]), .B1(\mx/mem[2][7] ), .B2(
        n2060), .ZN(n2161) );
  OAI22_X1 U2217 ( .A1(n2061), .A2(s_data_in_x[8]), .B1(\mx/mem[2][8] ), .B2(
        n2060), .ZN(n2162) );
  OAI22_X1 U2218 ( .A1(n2061), .A2(s_data_in_x[9]), .B1(\mx/mem[2][9] ), .B2(
        n2060), .ZN(n2163) );
  OAI22_X1 U2219 ( .A1(n2061), .A2(s_data_in_x[10]), .B1(\mx/mem[2][10] ), 
        .B2(n2060), .ZN(n2164) );
  OAI22_X1 U2220 ( .A1(n2061), .A2(s_data_in_x[11]), .B1(\mx/mem[2][11] ), 
        .B2(n2060), .ZN(n2165) );
  OAI22_X1 U2221 ( .A1(n2061), .A2(s_data_in_x[12]), .B1(\mx/mem[2][12] ), 
        .B2(n2060), .ZN(n2166) );
  OAI22_X1 U2222 ( .A1(n2061), .A2(s_data_in_x[13]), .B1(\mx/mem[2][13] ), 
        .B2(n2060), .ZN(n2167) );
  OAI22_X1 U2223 ( .A1(n2061), .A2(s_data_in_x[14]), .B1(\mx/mem[2][14] ), 
        .B2(n2060), .ZN(n2168) );
  OAI22_X1 U2224 ( .A1(n2061), .A2(s_data_in_x[15]), .B1(\mx/mem[2][15] ), 
        .B2(n2060), .ZN(n2169) );
  NOR2_X2 U2225 ( .A1(n2082), .A2(n2071), .ZN(n2062) );
  OAI22_X1 U2226 ( .A1(n2063), .A2(s_data_in_x[0]), .B1(\mx/mem[3][0] ), .B2(
        n2062), .ZN(n2170) );
  OAI22_X1 U2227 ( .A1(n2063), .A2(s_data_in_x[1]), .B1(\mx/mem[3][1] ), .B2(
        n2062), .ZN(n2171) );
  OAI22_X1 U2228 ( .A1(n2063), .A2(s_data_in_x[2]), .B1(\mx/mem[3][2] ), .B2(
        n2062), .ZN(n2172) );
  OAI22_X1 U2229 ( .A1(n2063), .A2(s_data_in_x[3]), .B1(\mx/mem[3][3] ), .B2(
        n2062), .ZN(n2173) );
  OAI22_X1 U2230 ( .A1(n2063), .A2(s_data_in_x[4]), .B1(\mx/mem[3][4] ), .B2(
        n2062), .ZN(n2174) );
  OAI22_X1 U2231 ( .A1(n2063), .A2(s_data_in_x[5]), .B1(\mx/mem[3][5] ), .B2(
        n2062), .ZN(n2175) );
  OAI22_X1 U2232 ( .A1(n2063), .A2(s_data_in_x[6]), .B1(\mx/mem[3][6] ), .B2(
        n2062), .ZN(n2176) );
  OAI22_X1 U2233 ( .A1(n2063), .A2(s_data_in_x[7]), .B1(\mx/mem[3][7] ), .B2(
        n2062), .ZN(n2177) );
  OAI22_X1 U2234 ( .A1(n2063), .A2(s_data_in_x[8]), .B1(\mx/mem[3][8] ), .B2(
        n2062), .ZN(n2178) );
  OAI22_X1 U2235 ( .A1(n2063), .A2(s_data_in_x[9]), .B1(\mx/mem[3][9] ), .B2(
        n2062), .ZN(n2179) );
  OAI22_X1 U2236 ( .A1(n2063), .A2(s_data_in_x[10]), .B1(\mx/mem[3][10] ), 
        .B2(n2062), .ZN(n2180) );
  OAI22_X1 U2237 ( .A1(n2063), .A2(s_data_in_x[11]), .B1(\mx/mem[3][11] ), 
        .B2(n2062), .ZN(n2181) );
  OAI22_X1 U2238 ( .A1(n2063), .A2(s_data_in_x[12]), .B1(\mx/mem[3][12] ), 
        .B2(n2062), .ZN(n2182) );
  OAI22_X1 U2239 ( .A1(n2063), .A2(s_data_in_x[13]), .B1(\mx/mem[3][13] ), 
        .B2(n2062), .ZN(n2183) );
  OAI22_X1 U2240 ( .A1(n2063), .A2(s_data_in_x[14]), .B1(\mx/mem[3][14] ), 
        .B2(n2062), .ZN(n2184) );
  OAI22_X1 U2241 ( .A1(n2063), .A2(s_data_in_x[15]), .B1(\mx/mem[3][15] ), 
        .B2(n2062), .ZN(n2185) );
  NOR2_X2 U2242 ( .A1(n2087), .A2(n2068), .ZN(n2064) );
  OAI22_X1 U2243 ( .A1(n2065), .A2(s_data_in_x[0]), .B1(\mx/mem[4][0] ), .B2(
        n2064), .ZN(n2186) );
  OAI22_X1 U2244 ( .A1(n2065), .A2(s_data_in_x[1]), .B1(\mx/mem[4][1] ), .B2(
        n2064), .ZN(n2187) );
  OAI22_X1 U2245 ( .A1(n2065), .A2(s_data_in_x[2]), .B1(\mx/mem[4][2] ), .B2(
        n2064), .ZN(n2188) );
  OAI22_X1 U2246 ( .A1(n2065), .A2(s_data_in_x[3]), .B1(\mx/mem[4][3] ), .B2(
        n2064), .ZN(n2189) );
  OAI22_X1 U2247 ( .A1(n2065), .A2(s_data_in_x[4]), .B1(\mx/mem[4][4] ), .B2(
        n2064), .ZN(n2190) );
  OAI22_X1 U2248 ( .A1(n2065), .A2(s_data_in_x[5]), .B1(\mx/mem[4][5] ), .B2(
        n2064), .ZN(n2191) );
  OAI22_X1 U2249 ( .A1(n2065), .A2(s_data_in_x[6]), .B1(\mx/mem[4][6] ), .B2(
        n2064), .ZN(n2192) );
  OAI22_X1 U2250 ( .A1(n2065), .A2(s_data_in_x[7]), .B1(\mx/mem[4][7] ), .B2(
        n2064), .ZN(n2193) );
  OAI22_X1 U2251 ( .A1(n2065), .A2(s_data_in_x[8]), .B1(\mx/mem[4][8] ), .B2(
        n2064), .ZN(n2194) );
  OAI22_X1 U2252 ( .A1(n2065), .A2(s_data_in_x[9]), .B1(\mx/mem[4][9] ), .B2(
        n2064), .ZN(n2195) );
  OAI22_X1 U2253 ( .A1(n2065), .A2(s_data_in_x[10]), .B1(\mx/mem[4][10] ), 
        .B2(n2064), .ZN(n2196) );
  OAI22_X1 U2254 ( .A1(n2065), .A2(s_data_in_x[11]), .B1(\mx/mem[4][11] ), 
        .B2(n2064), .ZN(n2197) );
  OAI22_X1 U2255 ( .A1(n2065), .A2(s_data_in_x[12]), .B1(\mx/mem[4][12] ), 
        .B2(n2064), .ZN(n2198) );
  OAI22_X1 U2256 ( .A1(n2065), .A2(s_data_in_x[13]), .B1(\mx/mem[4][13] ), 
        .B2(n2064), .ZN(n2199) );
  OAI22_X1 U2257 ( .A1(n2065), .A2(s_data_in_x[14]), .B1(\mx/mem[4][14] ), 
        .B2(n2064), .ZN(n2200) );
  OAI22_X1 U2258 ( .A1(n2065), .A2(s_data_in_x[15]), .B1(\mx/mem[4][15] ), 
        .B2(n2064), .ZN(n2201) );
  NOR2_X2 U2259 ( .A1(n2087), .A2(n2071), .ZN(n2066) );
  OAI22_X1 U2260 ( .A1(n2067), .A2(s_data_in_x[0]), .B1(\mx/mem[5][0] ), .B2(
        n2066), .ZN(n2202) );
  OAI22_X1 U2261 ( .A1(n2067), .A2(s_data_in_x[1]), .B1(\mx/mem[5][1] ), .B2(
        n2066), .ZN(n2203) );
  OAI22_X1 U2262 ( .A1(n2067), .A2(s_data_in_x[2]), .B1(\mx/mem[5][2] ), .B2(
        n2066), .ZN(n2204) );
  OAI22_X1 U2263 ( .A1(n2067), .A2(s_data_in_x[3]), .B1(\mx/mem[5][3] ), .B2(
        n2066), .ZN(n2205) );
  OAI22_X1 U2264 ( .A1(n2067), .A2(s_data_in_x[4]), .B1(\mx/mem[5][4] ), .B2(
        n2066), .ZN(n2206) );
  OAI22_X1 U2265 ( .A1(n2067), .A2(s_data_in_x[5]), .B1(\mx/mem[5][5] ), .B2(
        n2066), .ZN(n2207) );
  OAI22_X1 U2266 ( .A1(n2067), .A2(s_data_in_x[6]), .B1(\mx/mem[5][6] ), .B2(
        n2066), .ZN(n2208) );
  OAI22_X1 U2267 ( .A1(n2067), .A2(s_data_in_x[7]), .B1(\mx/mem[5][7] ), .B2(
        n2066), .ZN(n2209) );
  OAI22_X1 U2268 ( .A1(n2067), .A2(s_data_in_x[8]), .B1(\mx/mem[5][8] ), .B2(
        n2066), .ZN(n2210) );
  OAI22_X1 U2269 ( .A1(n2067), .A2(s_data_in_x[9]), .B1(\mx/mem[5][9] ), .B2(
        n2066), .ZN(n2211) );
  OAI22_X1 U2270 ( .A1(n2067), .A2(s_data_in_x[10]), .B1(\mx/mem[5][10] ), 
        .B2(n2066), .ZN(n2212) );
  OAI22_X1 U2271 ( .A1(n2067), .A2(s_data_in_x[11]), .B1(\mx/mem[5][11] ), 
        .B2(n2066), .ZN(n2213) );
  OAI22_X1 U2272 ( .A1(n2067), .A2(s_data_in_x[12]), .B1(\mx/mem[5][12] ), 
        .B2(n2066), .ZN(n2214) );
  OAI22_X1 U2273 ( .A1(n2067), .A2(s_data_in_x[13]), .B1(\mx/mem[5][13] ), 
        .B2(n2066), .ZN(n2215) );
  OAI22_X1 U2274 ( .A1(n2067), .A2(s_data_in_x[14]), .B1(\mx/mem[5][14] ), 
        .B2(n2066), .ZN(n2216) );
  OAI22_X1 U2275 ( .A1(n2067), .A2(s_data_in_x[15]), .B1(\mx/mem[5][15] ), 
        .B2(n2066), .ZN(n2217) );
  NOR2_X2 U2276 ( .A1(n2094), .A2(n2068), .ZN(n2069) );
  OAI22_X1 U2277 ( .A1(n2070), .A2(s_data_in_x[0]), .B1(\mx/mem[6][0] ), .B2(
        n2069), .ZN(n2218) );
  OAI22_X1 U2278 ( .A1(n2070), .A2(s_data_in_x[1]), .B1(\mx/mem[6][1] ), .B2(
        n2069), .ZN(n2219) );
  OAI22_X1 U2279 ( .A1(n2070), .A2(s_data_in_x[2]), .B1(\mx/mem[6][2] ), .B2(
        n2069), .ZN(n2220) );
  OAI22_X1 U2280 ( .A1(n2070), .A2(s_data_in_x[3]), .B1(\mx/mem[6][3] ), .B2(
        n2069), .ZN(n2221) );
  OAI22_X1 U2281 ( .A1(n2070), .A2(s_data_in_x[4]), .B1(\mx/mem[6][4] ), .B2(
        n2069), .ZN(n2222) );
  OAI22_X1 U2282 ( .A1(n2070), .A2(s_data_in_x[5]), .B1(\mx/mem[6][5] ), .B2(
        n2069), .ZN(n2223) );
  OAI22_X1 U2283 ( .A1(n2070), .A2(s_data_in_x[6]), .B1(\mx/mem[6][6] ), .B2(
        n2069), .ZN(n2224) );
  OAI22_X1 U2284 ( .A1(n2070), .A2(s_data_in_x[7]), .B1(\mx/mem[6][7] ), .B2(
        n2069), .ZN(n2225) );
  OAI22_X1 U2285 ( .A1(n2070), .A2(s_data_in_x[8]), .B1(\mx/mem[6][8] ), .B2(
        n2069), .ZN(n2226) );
  OAI22_X1 U2286 ( .A1(n2070), .A2(s_data_in_x[9]), .B1(\mx/mem[6][9] ), .B2(
        n2069), .ZN(n2227) );
  OAI22_X1 U2287 ( .A1(n2070), .A2(s_data_in_x[10]), .B1(\mx/mem[6][10] ), 
        .B2(n2069), .ZN(n2228) );
  OAI22_X1 U2288 ( .A1(n2070), .A2(s_data_in_x[11]), .B1(\mx/mem[6][11] ), 
        .B2(n2069), .ZN(n2229) );
  OAI22_X1 U2289 ( .A1(n2070), .A2(s_data_in_x[12]), .B1(\mx/mem[6][12] ), 
        .B2(n2069), .ZN(n2230) );
  OAI22_X1 U2290 ( .A1(n2070), .A2(s_data_in_x[13]), .B1(\mx/mem[6][13] ), 
        .B2(n2069), .ZN(n2231) );
  OAI22_X1 U2291 ( .A1(n2070), .A2(s_data_in_x[14]), .B1(\mx/mem[6][14] ), 
        .B2(n2069), .ZN(n2232) );
  OAI22_X1 U2292 ( .A1(n2070), .A2(s_data_in_x[15]), .B1(\mx/mem[6][15] ), 
        .B2(n2069), .ZN(n2233) );
  NOR2_X2 U2293 ( .A1(n2094), .A2(n2071), .ZN(n2072) );
  OAI22_X1 U2294 ( .A1(n2073), .A2(s_data_in_x[0]), .B1(\mx/mem[7][0] ), .B2(
        n2072), .ZN(n2234) );
  OAI22_X1 U2295 ( .A1(n2073), .A2(s_data_in_x[1]), .B1(\mx/mem[7][1] ), .B2(
        n2072), .ZN(n2235) );
  OAI22_X1 U2296 ( .A1(n2073), .A2(s_data_in_x[2]), .B1(\mx/mem[7][2] ), .B2(
        n2072), .ZN(n2236) );
  OAI22_X1 U2297 ( .A1(n2073), .A2(s_data_in_x[3]), .B1(\mx/mem[7][3] ), .B2(
        n2072), .ZN(n2237) );
  OAI22_X1 U2298 ( .A1(n2073), .A2(s_data_in_x[4]), .B1(\mx/mem[7][4] ), .B2(
        n2072), .ZN(n2238) );
  OAI22_X1 U2299 ( .A1(n2073), .A2(s_data_in_x[5]), .B1(\mx/mem[7][5] ), .B2(
        n2072), .ZN(n2239) );
  OAI22_X1 U2300 ( .A1(n2073), .A2(s_data_in_x[6]), .B1(\mx/mem[7][6] ), .B2(
        n2072), .ZN(n2240) );
  OAI22_X1 U2301 ( .A1(n2073), .A2(s_data_in_x[7]), .B1(\mx/mem[7][7] ), .B2(
        n2072), .ZN(n2241) );
  OAI22_X1 U2302 ( .A1(n2073), .A2(s_data_in_x[8]), .B1(\mx/mem[7][8] ), .B2(
        n2072), .ZN(n2242) );
  OAI22_X1 U2303 ( .A1(n2073), .A2(s_data_in_x[9]), .B1(\mx/mem[7][9] ), .B2(
        n2072), .ZN(n2243) );
  OAI22_X1 U2304 ( .A1(n2073), .A2(s_data_in_x[10]), .B1(\mx/mem[7][10] ), 
        .B2(n2072), .ZN(n2244) );
  OAI22_X1 U2305 ( .A1(n2073), .A2(s_data_in_x[11]), .B1(\mx/mem[7][11] ), 
        .B2(n2072), .ZN(n2245) );
  OAI22_X1 U2306 ( .A1(n2073), .A2(s_data_in_x[12]), .B1(\mx/mem[7][12] ), 
        .B2(n2072), .ZN(n2246) );
  OAI22_X1 U2307 ( .A1(n2073), .A2(s_data_in_x[13]), .B1(\mx/mem[7][13] ), 
        .B2(n2072), .ZN(n2247) );
  OAI22_X1 U2308 ( .A1(n2073), .A2(s_data_in_x[14]), .B1(\mx/mem[7][14] ), 
        .B2(n2072), .ZN(n2248) );
  OAI22_X1 U2309 ( .A1(n2073), .A2(s_data_in_x[15]), .B1(\mx/mem[7][15] ), 
        .B2(n2072), .ZN(n2249) );
  NAND2_X1 U2310 ( .A1(n2076), .A2(n2108), .ZN(n2090) );
  NOR2_X2 U2311 ( .A1(n2077), .A2(n2090), .ZN(n2074) );
  OAI22_X1 U2312 ( .A1(n2075), .A2(s_data_in_x[0]), .B1(\mx/mem[8][0] ), .B2(
        n2074), .ZN(n2250) );
  OAI22_X1 U2313 ( .A1(n2075), .A2(s_data_in_x[1]), .B1(\mx/mem[8][1] ), .B2(
        n2074), .ZN(n2251) );
  OAI22_X1 U2314 ( .A1(n2075), .A2(s_data_in_x[2]), .B1(\mx/mem[8][2] ), .B2(
        n2074), .ZN(n2252) );
  OAI22_X1 U2315 ( .A1(n2075), .A2(s_data_in_x[3]), .B1(\mx/mem[8][3] ), .B2(
        n2074), .ZN(n2253) );
  OAI22_X1 U2316 ( .A1(n2075), .A2(s_data_in_x[4]), .B1(\mx/mem[8][4] ), .B2(
        n2074), .ZN(n2254) );
  OAI22_X1 U2317 ( .A1(n2075), .A2(s_data_in_x[5]), .B1(\mx/mem[8][5] ), .B2(
        n2074), .ZN(n2255) );
  OAI22_X1 U2318 ( .A1(n2075), .A2(s_data_in_x[6]), .B1(\mx/mem[8][6] ), .B2(
        n2074), .ZN(n2256) );
  OAI22_X1 U2319 ( .A1(n2075), .A2(s_data_in_x[7]), .B1(\mx/mem[8][7] ), .B2(
        n2074), .ZN(n2257) );
  OAI22_X1 U2320 ( .A1(n2075), .A2(s_data_in_x[8]), .B1(\mx/mem[8][8] ), .B2(
        n2074), .ZN(n2258) );
  OAI22_X1 U2321 ( .A1(n2075), .A2(s_data_in_x[9]), .B1(\mx/mem[8][9] ), .B2(
        n2074), .ZN(n2259) );
  OAI22_X1 U2322 ( .A1(n2075), .A2(s_data_in_x[10]), .B1(\mx/mem[8][10] ), 
        .B2(n2074), .ZN(n2260) );
  OAI22_X1 U2323 ( .A1(n2075), .A2(s_data_in_x[11]), .B1(\mx/mem[8][11] ), 
        .B2(n2074), .ZN(n2261) );
  OAI22_X1 U2324 ( .A1(n2075), .A2(s_data_in_x[12]), .B1(\mx/mem[8][12] ), 
        .B2(n2074), .ZN(n2262) );
  OAI22_X1 U2325 ( .A1(n2075), .A2(s_data_in_x[13]), .B1(\mx/mem[8][13] ), 
        .B2(n2074), .ZN(n2263) );
  OAI22_X1 U2326 ( .A1(n2075), .A2(s_data_in_x[14]), .B1(\mx/mem[8][14] ), 
        .B2(n2074), .ZN(n2264) );
  OAI22_X1 U2327 ( .A1(n2075), .A2(s_data_in_x[15]), .B1(\mx/mem[8][15] ), 
        .B2(n2074), .ZN(n2265) );
  NAND2_X1 U2328 ( .A1(n2076), .A2(w_write_addr_x[0]), .ZN(n2093) );
  NOR2_X2 U2329 ( .A1(n2077), .A2(n2093), .ZN(n2078) );
  OAI22_X1 U2330 ( .A1(n2079), .A2(s_data_in_x[0]), .B1(\mx/mem[9][0] ), .B2(
        n2078), .ZN(n2266) );
  OAI22_X1 U2331 ( .A1(n2079), .A2(s_data_in_x[1]), .B1(\mx/mem[9][1] ), .B2(
        n2078), .ZN(n2267) );
  OAI22_X1 U2332 ( .A1(n2079), .A2(s_data_in_x[2]), .B1(\mx/mem[9][2] ), .B2(
        n2078), .ZN(n2268) );
  OAI22_X1 U2333 ( .A1(n2079), .A2(s_data_in_x[3]), .B1(\mx/mem[9][3] ), .B2(
        n2078), .ZN(n2269) );
  OAI22_X1 U2334 ( .A1(n2079), .A2(s_data_in_x[4]), .B1(\mx/mem[9][4] ), .B2(
        n2078), .ZN(n2270) );
  OAI22_X1 U2335 ( .A1(n2079), .A2(s_data_in_x[5]), .B1(\mx/mem[9][5] ), .B2(
        n2078), .ZN(n2271) );
  OAI22_X1 U2336 ( .A1(n2079), .A2(s_data_in_x[6]), .B1(\mx/mem[9][6] ), .B2(
        n2078), .ZN(n2272) );
  OAI22_X1 U2337 ( .A1(n2079), .A2(s_data_in_x[7]), .B1(\mx/mem[9][7] ), .B2(
        n2078), .ZN(n2273) );
  OAI22_X1 U2338 ( .A1(n2079), .A2(s_data_in_x[8]), .B1(\mx/mem[9][8] ), .B2(
        n2078), .ZN(n2274) );
  OAI22_X1 U2339 ( .A1(n2079), .A2(s_data_in_x[9]), .B1(\mx/mem[9][9] ), .B2(
        n2078), .ZN(n2275) );
  OAI22_X1 U2340 ( .A1(n2079), .A2(s_data_in_x[10]), .B1(\mx/mem[9][10] ), 
        .B2(n2078), .ZN(n2276) );
  OAI22_X1 U2341 ( .A1(n2079), .A2(s_data_in_x[11]), .B1(\mx/mem[9][11] ), 
        .B2(n2078), .ZN(n2277) );
  OAI22_X1 U2342 ( .A1(n2079), .A2(s_data_in_x[12]), .B1(\mx/mem[9][12] ), 
        .B2(n2078), .ZN(n2278) );
  OAI22_X1 U2343 ( .A1(n2079), .A2(s_data_in_x[13]), .B1(\mx/mem[9][13] ), 
        .B2(n2078), .ZN(n2279) );
  OAI22_X1 U2344 ( .A1(n2079), .A2(s_data_in_x[14]), .B1(\mx/mem[9][14] ), 
        .B2(n2078), .ZN(n2280) );
  OAI22_X1 U2345 ( .A1(n2079), .A2(s_data_in_x[15]), .B1(\mx/mem[9][15] ), 
        .B2(n2078), .ZN(n2281) );
  NOR2_X2 U2346 ( .A1(n2082), .A2(n2090), .ZN(n2080) );
  OAI22_X1 U2347 ( .A1(n2081), .A2(s_data_in_x[0]), .B1(\mx/mem[10][0] ), .B2(
        n2080), .ZN(n2282) );
  OAI22_X1 U2348 ( .A1(n2081), .A2(s_data_in_x[1]), .B1(\mx/mem[10][1] ), .B2(
        n2080), .ZN(n2283) );
  OAI22_X1 U2349 ( .A1(n2081), .A2(s_data_in_x[2]), .B1(\mx/mem[10][2] ), .B2(
        n2080), .ZN(n2284) );
  OAI22_X1 U2350 ( .A1(n2081), .A2(s_data_in_x[3]), .B1(\mx/mem[10][3] ), .B2(
        n2080), .ZN(n2285) );
  OAI22_X1 U2351 ( .A1(n2081), .A2(s_data_in_x[4]), .B1(\mx/mem[10][4] ), .B2(
        n2080), .ZN(n2286) );
  OAI22_X1 U2352 ( .A1(n2081), .A2(s_data_in_x[5]), .B1(\mx/mem[10][5] ), .B2(
        n2080), .ZN(n2287) );
  OAI22_X1 U2353 ( .A1(n2081), .A2(s_data_in_x[6]), .B1(\mx/mem[10][6] ), .B2(
        n2080), .ZN(n2288) );
  OAI22_X1 U2354 ( .A1(n2081), .A2(s_data_in_x[7]), .B1(\mx/mem[10][7] ), .B2(
        n2080), .ZN(n2289) );
  OAI22_X1 U2355 ( .A1(n2081), .A2(s_data_in_x[8]), .B1(\mx/mem[10][8] ), .B2(
        n2080), .ZN(n2290) );
  OAI22_X1 U2356 ( .A1(n2081), .A2(s_data_in_x[9]), .B1(\mx/mem[10][9] ), .B2(
        n2080), .ZN(n2291) );
  OAI22_X1 U2357 ( .A1(n2081), .A2(s_data_in_x[10]), .B1(\mx/mem[10][10] ), 
        .B2(n2080), .ZN(n2292) );
  OAI22_X1 U2358 ( .A1(n2081), .A2(s_data_in_x[11]), .B1(\mx/mem[10][11] ), 
        .B2(n2080), .ZN(n2293) );
  OAI22_X1 U2359 ( .A1(n2081), .A2(s_data_in_x[12]), .B1(\mx/mem[10][12] ), 
        .B2(n2080), .ZN(n2294) );
  OAI22_X1 U2360 ( .A1(n2081), .A2(s_data_in_x[13]), .B1(\mx/mem[10][13] ), 
        .B2(n2080), .ZN(n2295) );
  OAI22_X1 U2361 ( .A1(n2081), .A2(s_data_in_x[14]), .B1(\mx/mem[10][14] ), 
        .B2(n2080), .ZN(n2296) );
  OAI22_X1 U2362 ( .A1(n2081), .A2(s_data_in_x[15]), .B1(\mx/mem[10][15] ), 
        .B2(n2080), .ZN(n2297) );
  NOR2_X2 U2363 ( .A1(n2082), .A2(n2093), .ZN(n2083) );
  OAI22_X1 U2364 ( .A1(n2084), .A2(s_data_in_x[0]), .B1(\mx/mem[11][0] ), .B2(
        n2083), .ZN(n2298) );
  OAI22_X1 U2365 ( .A1(n2084), .A2(s_data_in_x[1]), .B1(\mx/mem[11][1] ), .B2(
        n2083), .ZN(n2299) );
  OAI22_X1 U2366 ( .A1(n2084), .A2(s_data_in_x[2]), .B1(\mx/mem[11][2] ), .B2(
        n2083), .ZN(n2300) );
  OAI22_X1 U2367 ( .A1(n2084), .A2(s_data_in_x[3]), .B1(\mx/mem[11][3] ), .B2(
        n2083), .ZN(n2301) );
  OAI22_X1 U2368 ( .A1(n2084), .A2(s_data_in_x[4]), .B1(\mx/mem[11][4] ), .B2(
        n2083), .ZN(n2302) );
  OAI22_X1 U2369 ( .A1(n2084), .A2(s_data_in_x[5]), .B1(\mx/mem[11][5] ), .B2(
        n2083), .ZN(n2303) );
  OAI22_X1 U2370 ( .A1(n2084), .A2(s_data_in_x[6]), .B1(\mx/mem[11][6] ), .B2(
        n2083), .ZN(n2304) );
  OAI22_X1 U2371 ( .A1(n2084), .A2(s_data_in_x[7]), .B1(\mx/mem[11][7] ), .B2(
        n2083), .ZN(n2305) );
  OAI22_X1 U2372 ( .A1(n2084), .A2(s_data_in_x[8]), .B1(\mx/mem[11][8] ), .B2(
        n2083), .ZN(n2306) );
  OAI22_X1 U2373 ( .A1(n2084), .A2(s_data_in_x[9]), .B1(\mx/mem[11][9] ), .B2(
        n2083), .ZN(n2307) );
  OAI22_X1 U2374 ( .A1(n2084), .A2(s_data_in_x[10]), .B1(\mx/mem[11][10] ), 
        .B2(n2083), .ZN(n2308) );
  OAI22_X1 U2375 ( .A1(n2084), .A2(s_data_in_x[11]), .B1(\mx/mem[11][11] ), 
        .B2(n2083), .ZN(n2309) );
  OAI22_X1 U2376 ( .A1(n2084), .A2(s_data_in_x[12]), .B1(\mx/mem[11][12] ), 
        .B2(n2083), .ZN(n2310) );
  OAI22_X1 U2377 ( .A1(n2084), .A2(s_data_in_x[13]), .B1(\mx/mem[11][13] ), 
        .B2(n2083), .ZN(n2311) );
  OAI22_X1 U2378 ( .A1(n2084), .A2(s_data_in_x[14]), .B1(\mx/mem[11][14] ), 
        .B2(n2083), .ZN(n2312) );
  OAI22_X1 U2379 ( .A1(n2084), .A2(s_data_in_x[15]), .B1(\mx/mem[11][15] ), 
        .B2(n2083), .ZN(n2313) );
  NOR2_X2 U2380 ( .A1(n2087), .A2(n2090), .ZN(n2085) );
  OAI22_X1 U2381 ( .A1(n2086), .A2(s_data_in_x[0]), .B1(\mx/mem[12][0] ), .B2(
        n2085), .ZN(n2314) );
  OAI22_X1 U2382 ( .A1(n2086), .A2(s_data_in_x[1]), .B1(\mx/mem[12][1] ), .B2(
        n2085), .ZN(n2315) );
  OAI22_X1 U2383 ( .A1(n2086), .A2(s_data_in_x[2]), .B1(\mx/mem[12][2] ), .B2(
        n2085), .ZN(n2316) );
  OAI22_X1 U2384 ( .A1(n2086), .A2(s_data_in_x[3]), .B1(\mx/mem[12][3] ), .B2(
        n2085), .ZN(n2317) );
  OAI22_X1 U2385 ( .A1(n2086), .A2(s_data_in_x[4]), .B1(\mx/mem[12][4] ), .B2(
        n2085), .ZN(n2318) );
  OAI22_X1 U2386 ( .A1(n2086), .A2(s_data_in_x[5]), .B1(\mx/mem[12][5] ), .B2(
        n2085), .ZN(n2319) );
  OAI22_X1 U2387 ( .A1(n2086), .A2(s_data_in_x[6]), .B1(\mx/mem[12][6] ), .B2(
        n2085), .ZN(n2320) );
  OAI22_X1 U2388 ( .A1(n2086), .A2(s_data_in_x[7]), .B1(\mx/mem[12][7] ), .B2(
        n2085), .ZN(n2321) );
  OAI22_X1 U2389 ( .A1(n2086), .A2(s_data_in_x[8]), .B1(\mx/mem[12][8] ), .B2(
        n2085), .ZN(n2322) );
  OAI22_X1 U2390 ( .A1(n2086), .A2(s_data_in_x[9]), .B1(\mx/mem[12][9] ), .B2(
        n2085), .ZN(n2323) );
  OAI22_X1 U2391 ( .A1(n2086), .A2(s_data_in_x[10]), .B1(\mx/mem[12][10] ), 
        .B2(n2085), .ZN(n2324) );
  OAI22_X1 U2392 ( .A1(n2086), .A2(s_data_in_x[11]), .B1(\mx/mem[12][11] ), 
        .B2(n2085), .ZN(n2325) );
  OAI22_X1 U2393 ( .A1(n2086), .A2(s_data_in_x[12]), .B1(\mx/mem[12][12] ), 
        .B2(n2085), .ZN(n2326) );
  OAI22_X1 U2394 ( .A1(n2086), .A2(s_data_in_x[13]), .B1(\mx/mem[12][13] ), 
        .B2(n2085), .ZN(n2327) );
  OAI22_X1 U2395 ( .A1(n2086), .A2(s_data_in_x[14]), .B1(\mx/mem[12][14] ), 
        .B2(n2085), .ZN(n2328) );
  OAI22_X1 U2396 ( .A1(n2086), .A2(s_data_in_x[15]), .B1(\mx/mem[12][15] ), 
        .B2(n2085), .ZN(n2329) );
  NOR2_X2 U2397 ( .A1(n2087), .A2(n2093), .ZN(n2088) );
  OAI22_X1 U2398 ( .A1(n2089), .A2(s_data_in_x[0]), .B1(\mx/mem[13][0] ), .B2(
        n2088), .ZN(n2330) );
  OAI22_X1 U2399 ( .A1(n2089), .A2(s_data_in_x[1]), .B1(\mx/mem[13][1] ), .B2(
        n2088), .ZN(n2331) );
  OAI22_X1 U2400 ( .A1(n2089), .A2(s_data_in_x[2]), .B1(\mx/mem[13][2] ), .B2(
        n2088), .ZN(n2332) );
  OAI22_X1 U2401 ( .A1(n2089), .A2(s_data_in_x[3]), .B1(\mx/mem[13][3] ), .B2(
        n2088), .ZN(n2333) );
  OAI22_X1 U2402 ( .A1(n2089), .A2(s_data_in_x[4]), .B1(\mx/mem[13][4] ), .B2(
        n2088), .ZN(n2334) );
  OAI22_X1 U2403 ( .A1(n2089), .A2(s_data_in_x[5]), .B1(\mx/mem[13][5] ), .B2(
        n2088), .ZN(n2335) );
  OAI22_X1 U2404 ( .A1(n2089), .A2(s_data_in_x[6]), .B1(\mx/mem[13][6] ), .B2(
        n2088), .ZN(n2336) );
  OAI22_X1 U2405 ( .A1(n2089), .A2(s_data_in_x[7]), .B1(\mx/mem[13][7] ), .B2(
        n2088), .ZN(n2337) );
  OAI22_X1 U2406 ( .A1(n2089), .A2(s_data_in_x[8]), .B1(\mx/mem[13][8] ), .B2(
        n2088), .ZN(n2338) );
  OAI22_X1 U2407 ( .A1(n2089), .A2(s_data_in_x[9]), .B1(\mx/mem[13][9] ), .B2(
        n2088), .ZN(n2339) );
  OAI22_X1 U2408 ( .A1(n2089), .A2(s_data_in_x[10]), .B1(\mx/mem[13][10] ), 
        .B2(n2088), .ZN(n2340) );
  OAI22_X1 U2409 ( .A1(n2089), .A2(s_data_in_x[11]), .B1(\mx/mem[13][11] ), 
        .B2(n2088), .ZN(n2341) );
  OAI22_X1 U2410 ( .A1(n2089), .A2(s_data_in_x[12]), .B1(\mx/mem[13][12] ), 
        .B2(n2088), .ZN(n2342) );
  OAI22_X1 U2411 ( .A1(n2089), .A2(s_data_in_x[13]), .B1(\mx/mem[13][13] ), 
        .B2(n2088), .ZN(n2343) );
  OAI22_X1 U2412 ( .A1(n2089), .A2(s_data_in_x[14]), .B1(\mx/mem[13][14] ), 
        .B2(n2088), .ZN(n2344) );
  OAI22_X1 U2413 ( .A1(n2089), .A2(s_data_in_x[15]), .B1(\mx/mem[13][15] ), 
        .B2(n2088), .ZN(n2345) );
  NOR2_X2 U2414 ( .A1(n2094), .A2(n2090), .ZN(n2091) );
  OAI22_X1 U2415 ( .A1(n2092), .A2(s_data_in_x[0]), .B1(\mx/mem[14][0] ), .B2(
        n2091), .ZN(n2346) );
  OAI22_X1 U2416 ( .A1(n2092), .A2(s_data_in_x[1]), .B1(\mx/mem[14][1] ), .B2(
        n2091), .ZN(n2347) );
  OAI22_X1 U2417 ( .A1(n2092), .A2(s_data_in_x[2]), .B1(\mx/mem[14][2] ), .B2(
        n2091), .ZN(n2348) );
  OAI22_X1 U2418 ( .A1(n2092), .A2(s_data_in_x[3]), .B1(\mx/mem[14][3] ), .B2(
        n2091), .ZN(n2349) );
  OAI22_X1 U2419 ( .A1(n2092), .A2(s_data_in_x[4]), .B1(\mx/mem[14][4] ), .B2(
        n2091), .ZN(n2350) );
  OAI22_X1 U2420 ( .A1(n2092), .A2(s_data_in_x[5]), .B1(\mx/mem[14][5] ), .B2(
        n2091), .ZN(n2351) );
  OAI22_X1 U2421 ( .A1(n2092), .A2(s_data_in_x[6]), .B1(\mx/mem[14][6] ), .B2(
        n2091), .ZN(n2352) );
  OAI22_X1 U2422 ( .A1(n2092), .A2(s_data_in_x[7]), .B1(\mx/mem[14][7] ), .B2(
        n2091), .ZN(n2353) );
  OAI22_X1 U2423 ( .A1(n2092), .A2(s_data_in_x[8]), .B1(\mx/mem[14][8] ), .B2(
        n2091), .ZN(n2354) );
  OAI22_X1 U2424 ( .A1(n2092), .A2(s_data_in_x[9]), .B1(\mx/mem[14][9] ), .B2(
        n2091), .ZN(n2355) );
  OAI22_X1 U2425 ( .A1(n2092), .A2(s_data_in_x[10]), .B1(\mx/mem[14][10] ), 
        .B2(n2091), .ZN(n2356) );
  OAI22_X1 U2426 ( .A1(n2092), .A2(s_data_in_x[11]), .B1(\mx/mem[14][11] ), 
        .B2(n2091), .ZN(n2357) );
  OAI22_X1 U2427 ( .A1(n2092), .A2(s_data_in_x[12]), .B1(\mx/mem[14][12] ), 
        .B2(n2091), .ZN(n2358) );
  OAI22_X1 U2428 ( .A1(n2092), .A2(s_data_in_x[13]), .B1(\mx/mem[14][13] ), 
        .B2(n2091), .ZN(n2359) );
  OAI22_X1 U2429 ( .A1(n2092), .A2(s_data_in_x[14]), .B1(\mx/mem[14][14] ), 
        .B2(n2091), .ZN(n2360) );
  OAI22_X1 U2430 ( .A1(n2092), .A2(s_data_in_x[15]), .B1(\mx/mem[14][15] ), 
        .B2(n2091), .ZN(n2361) );
  NOR2_X2 U2431 ( .A1(n2094), .A2(n2093), .ZN(n2095) );
  OAI22_X1 U2432 ( .A1(n2096), .A2(s_data_in_x[0]), .B1(\mx/mem[15][0] ), .B2(
        n2095), .ZN(n2362) );
  OAI22_X1 U2433 ( .A1(n2096), .A2(s_data_in_x[1]), .B1(\mx/mem[15][1] ), .B2(
        n2095), .ZN(n2363) );
  OAI22_X1 U2434 ( .A1(n2096), .A2(s_data_in_x[2]), .B1(\mx/mem[15][2] ), .B2(
        n2095), .ZN(n2364) );
  OAI22_X1 U2435 ( .A1(n2096), .A2(s_data_in_x[3]), .B1(\mx/mem[15][3] ), .B2(
        n2095), .ZN(n2365) );
  OAI22_X1 U2436 ( .A1(n2096), .A2(s_data_in_x[4]), .B1(\mx/mem[15][4] ), .B2(
        n2095), .ZN(n2366) );
  OAI22_X1 U2437 ( .A1(n2096), .A2(s_data_in_x[5]), .B1(\mx/mem[15][5] ), .B2(
        n2095), .ZN(n2367) );
  OAI22_X1 U2438 ( .A1(n2096), .A2(s_data_in_x[6]), .B1(\mx/mem[15][6] ), .B2(
        n2095), .ZN(n2368) );
  OAI22_X1 U2439 ( .A1(n2096), .A2(s_data_in_x[7]), .B1(\mx/mem[15][7] ), .B2(
        n2095), .ZN(n2369) );
  OAI22_X1 U2440 ( .A1(n2096), .A2(s_data_in_x[8]), .B1(\mx/mem[15][8] ), .B2(
        n2095), .ZN(n2370) );
  OAI22_X1 U2441 ( .A1(n2096), .A2(s_data_in_x[9]), .B1(\mx/mem[15][9] ), .B2(
        n2095), .ZN(n2371) );
  OAI22_X1 U2442 ( .A1(n2096), .A2(s_data_in_x[10]), .B1(\mx/mem[15][10] ), 
        .B2(n2095), .ZN(n2372) );
  OAI22_X1 U2443 ( .A1(n2096), .A2(s_data_in_x[11]), .B1(\mx/mem[15][11] ), 
        .B2(n2095), .ZN(n2373) );
  OAI22_X1 U2444 ( .A1(n2096), .A2(s_data_in_x[12]), .B1(\mx/mem[15][12] ), 
        .B2(n2095), .ZN(n2374) );
  OAI22_X1 U2445 ( .A1(n2096), .A2(s_data_in_x[13]), .B1(\mx/mem[15][13] ), 
        .B2(n2095), .ZN(n2375) );
  OAI22_X1 U2446 ( .A1(n2096), .A2(s_data_in_x[14]), .B1(\mx/mem[15][14] ), 
        .B2(n2095), .ZN(n2376) );
  OAI22_X1 U2447 ( .A1(n2096), .A2(s_data_in_x[15]), .B1(\mx/mem[15][15] ), 
        .B2(n2095), .ZN(n2377) );
endmodule

